// external module bram_r1_w1

// external module reg_r0_w1

// external module reg_r0_w1

// external module reg_r0_w1

// external module mult

