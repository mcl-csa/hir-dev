module kernel(	// matmul/matmul-hw.mlir:7651:3
  input  [15:0][31:0]  A_p0_rd_data,
  input  [255:0][31:0] B_p0_rd_data,
  input                t, clk, rst,
  output [15:0]        A_p0_addr_en,
  output [15:0][3:0]   A_p0_addr_data,
  output [15:0]        A_p0_rd_en,
  output [255:0]       B_p0_rd_en,
  output [15:0]        C_p0_addr_en,
  output [15:0][3:0]   C_p0_addr_data,
  output [15:0]        C_p0_wr_en,
  output [15:0][31:0]  C_p0_wr_data);

  wire [31:0]     _T;	// matmul/matmul-hw.mlir:23582:13
  wire            _T_0;	// matmul/matmul-hw.mlir:23581:13
  wire [3:0]      _T_1;	// matmul/matmul-hw.mlir:23580:13
  wire            _T_2;	// matmul/matmul-hw.mlir:23579:13
  wire            _T_3;	// matmul/matmul-hw.mlir:23563:13
  wire [31:0]     _T_4;	// matmul/matmul-hw.mlir:23539:13
  wire            _T_5;	// matmul/matmul-hw.mlir:23538:13
  wire            _T_6;	// matmul/matmul-hw.mlir:23521:13
  wire            _T_7;	// matmul/matmul-hw.mlir:23519:13
  wire            _T_8;	// matmul/matmul-hw.mlir:23518:13
  wire [31:0]     _T_9;	// matmul/matmul-hw.mlir:23509:13
  wire            _T_10;	// matmul/matmul-hw.mlir:23508:13
  wire            _T_11;	// matmul/matmul-hw.mlir:23491:13
  wire            _T_12;	// matmul/matmul-hw.mlir:23489:13
  wire            _T_13;	// matmul/matmul-hw.mlir:23488:13
  wire [31:0]     _T_14;	// matmul/matmul-hw.mlir:23479:13
  wire            _T_15;	// matmul/matmul-hw.mlir:23478:13
  wire            _T_16;	// matmul/matmul-hw.mlir:23461:13
  wire            _T_17;	// matmul/matmul-hw.mlir:23459:13
  wire            _T_18;	// matmul/matmul-hw.mlir:23458:13
  wire [31:0]     _T_19;	// matmul/matmul-hw.mlir:23449:13
  wire            _T_20;	// matmul/matmul-hw.mlir:23448:13
  wire            _T_21;	// matmul/matmul-hw.mlir:23431:13
  wire            _T_22;	// matmul/matmul-hw.mlir:23429:13
  wire            _T_23;	// matmul/matmul-hw.mlir:23428:13
  wire [31:0]     _T_24;	// matmul/matmul-hw.mlir:23419:13
  wire            _T_25;	// matmul/matmul-hw.mlir:23418:13
  wire            _T_26;	// matmul/matmul-hw.mlir:23401:13
  wire            _T_27;	// matmul/matmul-hw.mlir:23399:13
  wire            _T_28;	// matmul/matmul-hw.mlir:23398:13
  wire [31:0]     _T_29;	// matmul/matmul-hw.mlir:23389:13
  wire            _T_30;	// matmul/matmul-hw.mlir:23388:13
  wire            _T_31;	// matmul/matmul-hw.mlir:23371:13
  wire            _T_32;	// matmul/matmul-hw.mlir:23369:13
  wire            _T_33;	// matmul/matmul-hw.mlir:23368:13
  wire [31:0]     _T_34;	// matmul/matmul-hw.mlir:23359:13
  wire            _T_35;	// matmul/matmul-hw.mlir:23358:13
  wire            _T_36;	// matmul/matmul-hw.mlir:23341:13
  wire            _T_37;	// matmul/matmul-hw.mlir:23339:13
  wire            _T_38;	// matmul/matmul-hw.mlir:23338:13
  wire [31:0]     _T_39;	// matmul/matmul-hw.mlir:23329:13
  wire            _T_40;	// matmul/matmul-hw.mlir:23328:13
  wire            _T_41;	// matmul/matmul-hw.mlir:23311:13
  wire            _T_42;	// matmul/matmul-hw.mlir:23309:13
  wire            _T_43;	// matmul/matmul-hw.mlir:23308:13
  wire [31:0]     _T_44;	// matmul/matmul-hw.mlir:23299:13
  wire            _T_45;	// matmul/matmul-hw.mlir:23298:13
  wire            _T_46;	// matmul/matmul-hw.mlir:23281:13
  wire            _T_47;	// matmul/matmul-hw.mlir:23279:13
  wire            _T_48;	// matmul/matmul-hw.mlir:23278:13
  wire [31:0]     _T_49;	// matmul/matmul-hw.mlir:23269:13
  wire            _T_50;	// matmul/matmul-hw.mlir:23268:13
  wire            _T_51;	// matmul/matmul-hw.mlir:23251:13
  wire            _T_52;	// matmul/matmul-hw.mlir:23249:13
  wire            _T_53;	// matmul/matmul-hw.mlir:23248:13
  wire [31:0]     _T_54;	// matmul/matmul-hw.mlir:23239:13
  wire            _T_55;	// matmul/matmul-hw.mlir:23238:13
  wire            _T_56;	// matmul/matmul-hw.mlir:23221:13
  wire            _T_57;	// matmul/matmul-hw.mlir:23219:13
  wire            _T_58;	// matmul/matmul-hw.mlir:23218:13
  wire [31:0]     _T_59;	// matmul/matmul-hw.mlir:23209:13
  wire            _T_60;	// matmul/matmul-hw.mlir:23208:13
  wire            _T_61;	// matmul/matmul-hw.mlir:23191:13
  wire            _T_62;	// matmul/matmul-hw.mlir:23189:13
  wire            _T_63;	// matmul/matmul-hw.mlir:23188:13
  wire [31:0]     _T_64;	// matmul/matmul-hw.mlir:23179:13
  wire            _T_65;	// matmul/matmul-hw.mlir:23178:13
  wire            _T_66;	// matmul/matmul-hw.mlir:23161:13
  wire            _T_67;	// matmul/matmul-hw.mlir:23159:13
  wire            _T_68;	// matmul/matmul-hw.mlir:23158:13
  wire [31:0]     _T_69;	// matmul/matmul-hw.mlir:23149:13
  wire            _T_70;	// matmul/matmul-hw.mlir:23148:13
  wire            _T_71;	// matmul/matmul-hw.mlir:23131:13
  wire            _T_72;	// matmul/matmul-hw.mlir:23129:13
  wire            _T_73;	// matmul/matmul-hw.mlir:23128:13
  wire [31:0]     _T_74;	// matmul/matmul-hw.mlir:23119:13
  wire            _T_75;	// matmul/matmul-hw.mlir:23118:13
  wire            _T_76;	// matmul/matmul-hw.mlir:23101:13
  wire            _T_77;	// matmul/matmul-hw.mlir:23099:13
  wire            _T_78;	// matmul/matmul-hw.mlir:23098:13
  wire [31:0]     _T_79;	// matmul/matmul-hw.mlir:23089:13
  wire            _T_80;	// matmul/matmul-hw.mlir:23088:13
  wire            _T_81;	// matmul/matmul-hw.mlir:23071:13
  wire            _T_82;	// matmul/matmul-hw.mlir:23069:13
  wire            _T_83;	// matmul/matmul-hw.mlir:23068:13
  wire [31:0]     _T_84;	// matmul/matmul-hw.mlir:23067:13
  wire            _T_85;	// matmul/matmul-hw.mlir:23066:13
  wire [31:0]     _T_86;	// matmul/matmul-hw.mlir:22972:13
  wire            _T_87;	// matmul/matmul-hw.mlir:22971:13
  wire [3:0]      _T_88;	// matmul/matmul-hw.mlir:22970:13
  wire            _T_89;	// matmul/matmul-hw.mlir:22969:13
  wire            _T_90;	// matmul/matmul-hw.mlir:22953:13
  wire [31:0]     _T_91;	// matmul/matmul-hw.mlir:22929:13
  wire            _T_92;	// matmul/matmul-hw.mlir:22928:13
  wire            _T_93;	// matmul/matmul-hw.mlir:22911:13
  wire            _T_94;	// matmul/matmul-hw.mlir:22909:13
  wire            _T_95;	// matmul/matmul-hw.mlir:22908:13
  wire [31:0]     _T_96;	// matmul/matmul-hw.mlir:22899:13
  wire            _T_97;	// matmul/matmul-hw.mlir:22898:13
  wire            _T_98;	// matmul/matmul-hw.mlir:22881:13
  wire            _T_99;	// matmul/matmul-hw.mlir:22879:13
  wire            _T_100;	// matmul/matmul-hw.mlir:22878:13
  wire [31:0]     _T_101;	// matmul/matmul-hw.mlir:22869:13
  wire            _T_102;	// matmul/matmul-hw.mlir:22868:13
  wire            _T_103;	// matmul/matmul-hw.mlir:22851:13
  wire            _T_104;	// matmul/matmul-hw.mlir:22849:13
  wire            _T_105;	// matmul/matmul-hw.mlir:22848:13
  wire [31:0]     _T_106;	// matmul/matmul-hw.mlir:22839:13
  wire            _T_107;	// matmul/matmul-hw.mlir:22838:13
  wire            _T_108;	// matmul/matmul-hw.mlir:22821:13
  wire            _T_109;	// matmul/matmul-hw.mlir:22819:13
  wire            _T_110;	// matmul/matmul-hw.mlir:22818:13
  wire [31:0]     _T_111;	// matmul/matmul-hw.mlir:22809:13
  wire            _T_112;	// matmul/matmul-hw.mlir:22808:13
  wire            _T_113;	// matmul/matmul-hw.mlir:22791:13
  wire            _T_114;	// matmul/matmul-hw.mlir:22789:13
  wire            _T_115;	// matmul/matmul-hw.mlir:22788:13
  wire [31:0]     _T_116;	// matmul/matmul-hw.mlir:22779:13
  wire            _T_117;	// matmul/matmul-hw.mlir:22778:13
  wire            _T_118;	// matmul/matmul-hw.mlir:22761:13
  wire            _T_119;	// matmul/matmul-hw.mlir:22759:13
  wire            _T_120;	// matmul/matmul-hw.mlir:22758:13
  wire [31:0]     _T_121;	// matmul/matmul-hw.mlir:22749:13
  wire            _T_122;	// matmul/matmul-hw.mlir:22748:13
  wire            _T_123;	// matmul/matmul-hw.mlir:22731:13
  wire            _T_124;	// matmul/matmul-hw.mlir:22729:13
  wire            _T_125;	// matmul/matmul-hw.mlir:22728:13
  wire [31:0]     _T_126;	// matmul/matmul-hw.mlir:22719:13
  wire            _T_127;	// matmul/matmul-hw.mlir:22718:13
  wire            _T_128;	// matmul/matmul-hw.mlir:22701:13
  wire            _T_129;	// matmul/matmul-hw.mlir:22699:13
  wire            _T_130;	// matmul/matmul-hw.mlir:22698:13
  wire [31:0]     _T_131;	// matmul/matmul-hw.mlir:22689:13
  wire            _T_132;	// matmul/matmul-hw.mlir:22688:13
  wire            _T_133;	// matmul/matmul-hw.mlir:22671:13
  wire            _T_134;	// matmul/matmul-hw.mlir:22669:13
  wire            _T_135;	// matmul/matmul-hw.mlir:22668:13
  wire [31:0]     _T_136;	// matmul/matmul-hw.mlir:22659:13
  wire            _T_137;	// matmul/matmul-hw.mlir:22658:13
  wire            _T_138;	// matmul/matmul-hw.mlir:22641:13
  wire            _T_139;	// matmul/matmul-hw.mlir:22639:13
  wire            _T_140;	// matmul/matmul-hw.mlir:22638:13
  wire [31:0]     _T_141;	// matmul/matmul-hw.mlir:22629:13
  wire            _T_142;	// matmul/matmul-hw.mlir:22628:13
  wire            _T_143;	// matmul/matmul-hw.mlir:22611:13
  wire            _T_144;	// matmul/matmul-hw.mlir:22609:13
  wire            _T_145;	// matmul/matmul-hw.mlir:22608:13
  wire [31:0]     _T_146;	// matmul/matmul-hw.mlir:22599:13
  wire            _T_147;	// matmul/matmul-hw.mlir:22598:13
  wire            _T_148;	// matmul/matmul-hw.mlir:22581:13
  wire            _T_149;	// matmul/matmul-hw.mlir:22579:13
  wire            _T_150;	// matmul/matmul-hw.mlir:22578:13
  wire [31:0]     _T_151;	// matmul/matmul-hw.mlir:22569:13
  wire            _T_152;	// matmul/matmul-hw.mlir:22568:13
  wire            _T_153;	// matmul/matmul-hw.mlir:22551:13
  wire            _T_154;	// matmul/matmul-hw.mlir:22549:13
  wire            _T_155;	// matmul/matmul-hw.mlir:22548:13
  wire [31:0]     _T_156;	// matmul/matmul-hw.mlir:22539:13
  wire            _T_157;	// matmul/matmul-hw.mlir:22538:13
  wire            _T_158;	// matmul/matmul-hw.mlir:22521:13
  wire            _T_159;	// matmul/matmul-hw.mlir:22519:13
  wire            _T_160;	// matmul/matmul-hw.mlir:22518:13
  wire [31:0]     _T_161;	// matmul/matmul-hw.mlir:22509:13
  wire            _T_162;	// matmul/matmul-hw.mlir:22508:13
  wire            _T_163;	// matmul/matmul-hw.mlir:22491:13
  wire            _T_164;	// matmul/matmul-hw.mlir:22489:13
  wire            _T_165;	// matmul/matmul-hw.mlir:22488:13
  wire [31:0]     _T_166;	// matmul/matmul-hw.mlir:22479:13
  wire            _T_167;	// matmul/matmul-hw.mlir:22478:13
  wire            _T_168;	// matmul/matmul-hw.mlir:22461:13
  wire            _T_169;	// matmul/matmul-hw.mlir:22459:13
  wire            _T_170;	// matmul/matmul-hw.mlir:22458:13
  wire [31:0]     _T_171;	// matmul/matmul-hw.mlir:22457:13
  wire            _T_172;	// matmul/matmul-hw.mlir:22456:13
  wire [31:0]     _T_173;	// matmul/matmul-hw.mlir:22362:13
  wire            _T_174;	// matmul/matmul-hw.mlir:22361:13
  wire [3:0]      _T_175;	// matmul/matmul-hw.mlir:22360:13
  wire            _T_176;	// matmul/matmul-hw.mlir:22359:13
  wire            _T_177;	// matmul/matmul-hw.mlir:22343:13
  wire [31:0]     _T_178;	// matmul/matmul-hw.mlir:22319:13
  wire            _T_179;	// matmul/matmul-hw.mlir:22318:13
  wire            _T_180;	// matmul/matmul-hw.mlir:22301:13
  wire            _T_181;	// matmul/matmul-hw.mlir:22299:13
  wire            _T_182;	// matmul/matmul-hw.mlir:22298:13
  wire [31:0]     _T_183;	// matmul/matmul-hw.mlir:22289:13
  wire            _T_184;	// matmul/matmul-hw.mlir:22288:13
  wire            _T_185;	// matmul/matmul-hw.mlir:22271:13
  wire            _T_186;	// matmul/matmul-hw.mlir:22269:13
  wire            _T_187;	// matmul/matmul-hw.mlir:22268:13
  wire [31:0]     _T_188;	// matmul/matmul-hw.mlir:22259:13
  wire            _T_189;	// matmul/matmul-hw.mlir:22258:13
  wire            _T_190;	// matmul/matmul-hw.mlir:22241:13
  wire            _T_191;	// matmul/matmul-hw.mlir:22239:13
  wire            _T_192;	// matmul/matmul-hw.mlir:22238:13
  wire [31:0]     _T_193;	// matmul/matmul-hw.mlir:22229:13
  wire            _T_194;	// matmul/matmul-hw.mlir:22228:13
  wire            _T_195;	// matmul/matmul-hw.mlir:22211:13
  wire            _T_196;	// matmul/matmul-hw.mlir:22209:13
  wire            _T_197;	// matmul/matmul-hw.mlir:22208:13
  wire [31:0]     _T_198;	// matmul/matmul-hw.mlir:22199:13
  wire            _T_199;	// matmul/matmul-hw.mlir:22198:13
  wire            _T_200;	// matmul/matmul-hw.mlir:22181:13
  wire            _T_201;	// matmul/matmul-hw.mlir:22179:13
  wire            _T_202;	// matmul/matmul-hw.mlir:22178:13
  wire [31:0]     _T_203;	// matmul/matmul-hw.mlir:22169:13
  wire            _T_204;	// matmul/matmul-hw.mlir:22168:13
  wire            _T_205;	// matmul/matmul-hw.mlir:22151:13
  wire            _T_206;	// matmul/matmul-hw.mlir:22149:13
  wire            _T_207;	// matmul/matmul-hw.mlir:22148:13
  wire [31:0]     _T_208;	// matmul/matmul-hw.mlir:22139:13
  wire            _T_209;	// matmul/matmul-hw.mlir:22138:13
  wire            _T_210;	// matmul/matmul-hw.mlir:22121:13
  wire            _T_211;	// matmul/matmul-hw.mlir:22119:13
  wire            _T_212;	// matmul/matmul-hw.mlir:22118:13
  wire [31:0]     _T_213;	// matmul/matmul-hw.mlir:22109:13
  wire            _T_214;	// matmul/matmul-hw.mlir:22108:13
  wire            _T_215;	// matmul/matmul-hw.mlir:22091:13
  wire            _T_216;	// matmul/matmul-hw.mlir:22089:13
  wire            _T_217;	// matmul/matmul-hw.mlir:22088:13
  wire [31:0]     _T_218;	// matmul/matmul-hw.mlir:22079:13
  wire            _T_219;	// matmul/matmul-hw.mlir:22078:13
  wire            _T_220;	// matmul/matmul-hw.mlir:22061:13
  wire            _T_221;	// matmul/matmul-hw.mlir:22059:13
  wire            _T_222;	// matmul/matmul-hw.mlir:22058:13
  wire [31:0]     _T_223;	// matmul/matmul-hw.mlir:22049:13
  wire            _T_224;	// matmul/matmul-hw.mlir:22048:13
  wire            _T_225;	// matmul/matmul-hw.mlir:22031:13
  wire            _T_226;	// matmul/matmul-hw.mlir:22029:13
  wire            _T_227;	// matmul/matmul-hw.mlir:22028:13
  wire [31:0]     _T_228;	// matmul/matmul-hw.mlir:22019:13
  wire            _T_229;	// matmul/matmul-hw.mlir:22018:13
  wire            _T_230;	// matmul/matmul-hw.mlir:22001:13
  wire            _T_231;	// matmul/matmul-hw.mlir:21999:13
  wire            _T_232;	// matmul/matmul-hw.mlir:21998:13
  wire [31:0]     _T_233;	// matmul/matmul-hw.mlir:21989:13
  wire            _T_234;	// matmul/matmul-hw.mlir:21988:13
  wire            _T_235;	// matmul/matmul-hw.mlir:21971:13
  wire            _T_236;	// matmul/matmul-hw.mlir:21969:13
  wire            _T_237;	// matmul/matmul-hw.mlir:21968:13
  wire [31:0]     _T_238;	// matmul/matmul-hw.mlir:21959:13
  wire            _T_239;	// matmul/matmul-hw.mlir:21958:13
  wire            _T_240;	// matmul/matmul-hw.mlir:21941:13
  wire            _T_241;	// matmul/matmul-hw.mlir:21939:13
  wire            _T_242;	// matmul/matmul-hw.mlir:21938:13
  wire [31:0]     _T_243;	// matmul/matmul-hw.mlir:21929:13
  wire            _T_244;	// matmul/matmul-hw.mlir:21928:13
  wire            _T_245;	// matmul/matmul-hw.mlir:21911:13
  wire            _T_246;	// matmul/matmul-hw.mlir:21909:13
  wire            _T_247;	// matmul/matmul-hw.mlir:21908:13
  wire [31:0]     _T_248;	// matmul/matmul-hw.mlir:21899:13
  wire            _T_249;	// matmul/matmul-hw.mlir:21898:13
  wire            _T_250;	// matmul/matmul-hw.mlir:21881:13
  wire            _T_251;	// matmul/matmul-hw.mlir:21879:13
  wire            _T_252;	// matmul/matmul-hw.mlir:21878:13
  wire [31:0]     _T_253;	// matmul/matmul-hw.mlir:21869:13
  wire            _T_254;	// matmul/matmul-hw.mlir:21868:13
  wire            _T_255;	// matmul/matmul-hw.mlir:21851:13
  wire            _T_256;	// matmul/matmul-hw.mlir:21849:13
  wire            _T_257;	// matmul/matmul-hw.mlir:21848:13
  wire [31:0]     _T_258;	// matmul/matmul-hw.mlir:21847:13
  wire            _T_259;	// matmul/matmul-hw.mlir:21846:13
  wire [31:0]     _T_260;	// matmul/matmul-hw.mlir:21752:13
  wire            _T_261;	// matmul/matmul-hw.mlir:21751:13
  wire [3:0]      _T_262;	// matmul/matmul-hw.mlir:21750:13
  wire            _T_263;	// matmul/matmul-hw.mlir:21749:13
  wire            _T_264;	// matmul/matmul-hw.mlir:21733:13
  wire [31:0]     _T_265;	// matmul/matmul-hw.mlir:21709:13
  wire            _T_266;	// matmul/matmul-hw.mlir:21708:13
  wire            _T_267;	// matmul/matmul-hw.mlir:21691:13
  wire            _T_268;	// matmul/matmul-hw.mlir:21689:13
  wire            _T_269;	// matmul/matmul-hw.mlir:21688:13
  wire [31:0]     _T_270;	// matmul/matmul-hw.mlir:21679:13
  wire            _T_271;	// matmul/matmul-hw.mlir:21678:13
  wire            _T_272;	// matmul/matmul-hw.mlir:21661:13
  wire            _T_273;	// matmul/matmul-hw.mlir:21659:13
  wire            _T_274;	// matmul/matmul-hw.mlir:21658:13
  wire [31:0]     _T_275;	// matmul/matmul-hw.mlir:21649:13
  wire            _T_276;	// matmul/matmul-hw.mlir:21648:13
  wire            _T_277;	// matmul/matmul-hw.mlir:21631:13
  wire            _T_278;	// matmul/matmul-hw.mlir:21629:13
  wire            _T_279;	// matmul/matmul-hw.mlir:21628:13
  wire [31:0]     _T_280;	// matmul/matmul-hw.mlir:21619:13
  wire            _T_281;	// matmul/matmul-hw.mlir:21618:13
  wire            _T_282;	// matmul/matmul-hw.mlir:21601:13
  wire            _T_283;	// matmul/matmul-hw.mlir:21599:13
  wire            _T_284;	// matmul/matmul-hw.mlir:21598:13
  wire [31:0]     _T_285;	// matmul/matmul-hw.mlir:21589:13
  wire            _T_286;	// matmul/matmul-hw.mlir:21588:13
  wire            _T_287;	// matmul/matmul-hw.mlir:21571:13
  wire            _T_288;	// matmul/matmul-hw.mlir:21569:13
  wire            _T_289;	// matmul/matmul-hw.mlir:21568:13
  wire [31:0]     _T_290;	// matmul/matmul-hw.mlir:21559:13
  wire            _T_291;	// matmul/matmul-hw.mlir:21558:13
  wire            _T_292;	// matmul/matmul-hw.mlir:21541:13
  wire            _T_293;	// matmul/matmul-hw.mlir:21539:13
  wire            _T_294;	// matmul/matmul-hw.mlir:21538:13
  wire [31:0]     _T_295;	// matmul/matmul-hw.mlir:21529:13
  wire            _T_296;	// matmul/matmul-hw.mlir:21528:13
  wire            _T_297;	// matmul/matmul-hw.mlir:21511:13
  wire            _T_298;	// matmul/matmul-hw.mlir:21509:13
  wire            _T_299;	// matmul/matmul-hw.mlir:21508:13
  wire [31:0]     _T_300;	// matmul/matmul-hw.mlir:21499:13
  wire            _T_301;	// matmul/matmul-hw.mlir:21498:13
  wire            _T_302;	// matmul/matmul-hw.mlir:21481:13
  wire            _T_303;	// matmul/matmul-hw.mlir:21479:13
  wire            _T_304;	// matmul/matmul-hw.mlir:21478:13
  wire [31:0]     _T_305;	// matmul/matmul-hw.mlir:21469:13
  wire            _T_306;	// matmul/matmul-hw.mlir:21468:13
  wire            _T_307;	// matmul/matmul-hw.mlir:21451:13
  wire            _T_308;	// matmul/matmul-hw.mlir:21449:13
  wire            _T_309;	// matmul/matmul-hw.mlir:21448:13
  wire [31:0]     _T_310;	// matmul/matmul-hw.mlir:21439:13
  wire            _T_311;	// matmul/matmul-hw.mlir:21438:13
  wire            _T_312;	// matmul/matmul-hw.mlir:21421:13
  wire            _T_313;	// matmul/matmul-hw.mlir:21419:13
  wire            _T_314;	// matmul/matmul-hw.mlir:21418:13
  wire [31:0]     _T_315;	// matmul/matmul-hw.mlir:21409:13
  wire            _T_316;	// matmul/matmul-hw.mlir:21408:13
  wire            _T_317;	// matmul/matmul-hw.mlir:21391:13
  wire            _T_318;	// matmul/matmul-hw.mlir:21389:13
  wire            _T_319;	// matmul/matmul-hw.mlir:21388:13
  wire [31:0]     _T_320;	// matmul/matmul-hw.mlir:21379:13
  wire            _T_321;	// matmul/matmul-hw.mlir:21378:13
  wire            _T_322;	// matmul/matmul-hw.mlir:21361:13
  wire            _T_323;	// matmul/matmul-hw.mlir:21359:13
  wire            _T_324;	// matmul/matmul-hw.mlir:21358:13
  wire [31:0]     _T_325;	// matmul/matmul-hw.mlir:21349:13
  wire            _T_326;	// matmul/matmul-hw.mlir:21348:13
  wire            _T_327;	// matmul/matmul-hw.mlir:21331:13
  wire            _T_328;	// matmul/matmul-hw.mlir:21329:13
  wire            _T_329;	// matmul/matmul-hw.mlir:21328:13
  wire [31:0]     _T_330;	// matmul/matmul-hw.mlir:21319:13
  wire            _T_331;	// matmul/matmul-hw.mlir:21318:13
  wire            _T_332;	// matmul/matmul-hw.mlir:21301:13
  wire            _T_333;	// matmul/matmul-hw.mlir:21299:13
  wire            _T_334;	// matmul/matmul-hw.mlir:21298:13
  wire [31:0]     _T_335;	// matmul/matmul-hw.mlir:21289:13
  wire            _T_336;	// matmul/matmul-hw.mlir:21288:13
  wire            _T_337;	// matmul/matmul-hw.mlir:21271:13
  wire            _T_338;	// matmul/matmul-hw.mlir:21269:13
  wire            _T_339;	// matmul/matmul-hw.mlir:21268:13
  wire [31:0]     _T_340;	// matmul/matmul-hw.mlir:21259:13
  wire            _T_341;	// matmul/matmul-hw.mlir:21258:13
  wire            _T_342;	// matmul/matmul-hw.mlir:21241:13
  wire            _T_343;	// matmul/matmul-hw.mlir:21239:13
  wire            _T_344;	// matmul/matmul-hw.mlir:21238:13
  wire [31:0]     _T_345;	// matmul/matmul-hw.mlir:21237:13
  wire            _T_346;	// matmul/matmul-hw.mlir:21236:13
  wire [31:0]     _T_347;	// matmul/matmul-hw.mlir:21142:13
  wire            _T_348;	// matmul/matmul-hw.mlir:21141:13
  wire [3:0]      _T_349;	// matmul/matmul-hw.mlir:21140:13
  wire            _T_350;	// matmul/matmul-hw.mlir:21139:13
  wire            _T_351;	// matmul/matmul-hw.mlir:21123:13
  wire [31:0]     _T_352;	// matmul/matmul-hw.mlir:21114:13
  wire            _T_353;	// matmul/matmul-hw.mlir:21113:13
  wire            _T_354;	// matmul/matmul-hw.mlir:21096:13
  wire            _T_355;	// matmul/matmul-hw.mlir:21094:13
  wire            _T_356;	// matmul/matmul-hw.mlir:21093:13
  wire [31:0]     _T_357;	// matmul/matmul-hw.mlir:21084:13
  wire            _T_358;	// matmul/matmul-hw.mlir:21083:13
  wire            _T_359;	// matmul/matmul-hw.mlir:21066:13
  wire            _T_360;	// matmul/matmul-hw.mlir:21064:13
  wire            _T_361;	// matmul/matmul-hw.mlir:21063:13
  wire [31:0]     _T_362;	// matmul/matmul-hw.mlir:21054:13
  wire            _T_363;	// matmul/matmul-hw.mlir:21053:13
  wire            _T_364;	// matmul/matmul-hw.mlir:21036:13
  wire            _T_365;	// matmul/matmul-hw.mlir:21034:13
  wire            _T_366;	// matmul/matmul-hw.mlir:21033:13
  wire [31:0]     _T_367;	// matmul/matmul-hw.mlir:21024:13
  wire            _T_368;	// matmul/matmul-hw.mlir:21023:13
  wire            _T_369;	// matmul/matmul-hw.mlir:21006:13
  wire            _T_370;	// matmul/matmul-hw.mlir:21004:13
  wire            _T_371;	// matmul/matmul-hw.mlir:21003:13
  wire [31:0]     _T_372;	// matmul/matmul-hw.mlir:20994:13
  wire            _T_373;	// matmul/matmul-hw.mlir:20993:13
  wire            _T_374;	// matmul/matmul-hw.mlir:20976:13
  wire            _T_375;	// matmul/matmul-hw.mlir:20974:13
  wire            _T_376;	// matmul/matmul-hw.mlir:20973:13
  wire [31:0]     _T_377;	// matmul/matmul-hw.mlir:20964:13
  wire            _T_378;	// matmul/matmul-hw.mlir:20963:13
  wire            _T_379;	// matmul/matmul-hw.mlir:20946:13
  wire            _T_380;	// matmul/matmul-hw.mlir:20944:13
  wire            _T_381;	// matmul/matmul-hw.mlir:20943:13
  wire [31:0]     _T_382;	// matmul/matmul-hw.mlir:20934:13
  wire            _T_383;	// matmul/matmul-hw.mlir:20933:13
  wire            _T_384;	// matmul/matmul-hw.mlir:20916:13
  wire            _T_385;	// matmul/matmul-hw.mlir:20914:13
  wire            _T_386;	// matmul/matmul-hw.mlir:20913:13
  wire [31:0]     _T_387;	// matmul/matmul-hw.mlir:20904:13
  wire            _T_388;	// matmul/matmul-hw.mlir:20903:13
  wire            _T_389;	// matmul/matmul-hw.mlir:20886:13
  wire            _T_390;	// matmul/matmul-hw.mlir:20884:13
  wire            _T_391;	// matmul/matmul-hw.mlir:20883:13
  wire [31:0]     _T_392;	// matmul/matmul-hw.mlir:20874:13
  wire            _T_393;	// matmul/matmul-hw.mlir:20873:13
  wire            _T_394;	// matmul/matmul-hw.mlir:20856:13
  wire            _T_395;	// matmul/matmul-hw.mlir:20854:13
  wire            _T_396;	// matmul/matmul-hw.mlir:20853:13
  wire [31:0]     _T_397;	// matmul/matmul-hw.mlir:20844:13
  wire            _T_398;	// matmul/matmul-hw.mlir:20843:13
  wire            _T_399;	// matmul/matmul-hw.mlir:20826:13
  wire            _T_400;	// matmul/matmul-hw.mlir:20824:13
  wire            _T_401;	// matmul/matmul-hw.mlir:20823:13
  wire [31:0]     _T_402;	// matmul/matmul-hw.mlir:20814:13
  wire            _T_403;	// matmul/matmul-hw.mlir:20813:13
  wire            _T_404;	// matmul/matmul-hw.mlir:20796:13
  wire            _T_405;	// matmul/matmul-hw.mlir:20794:13
  wire            _T_406;	// matmul/matmul-hw.mlir:20793:13
  wire [31:0]     _T_407;	// matmul/matmul-hw.mlir:20784:13
  wire            _T_408;	// matmul/matmul-hw.mlir:20783:13
  wire            _T_409;	// matmul/matmul-hw.mlir:20766:13
  wire            _T_410;	// matmul/matmul-hw.mlir:20764:13
  wire            _T_411;	// matmul/matmul-hw.mlir:20763:13
  wire [31:0]     _T_412;	// matmul/matmul-hw.mlir:20754:13
  wire            _T_413;	// matmul/matmul-hw.mlir:20753:13
  wire            _T_414;	// matmul/matmul-hw.mlir:20736:13
  wire            _T_415;	// matmul/matmul-hw.mlir:20734:13
  wire            _T_416;	// matmul/matmul-hw.mlir:20733:13
  wire [31:0]     _T_417;	// matmul/matmul-hw.mlir:20724:13
  wire            _T_418;	// matmul/matmul-hw.mlir:20723:13
  wire            _T_419;	// matmul/matmul-hw.mlir:20706:13
  wire            _T_420;	// matmul/matmul-hw.mlir:20704:13
  wire            _T_421;	// matmul/matmul-hw.mlir:20703:13
  wire [31:0]     _T_422;	// matmul/matmul-hw.mlir:20694:13
  wire            _T_423;	// matmul/matmul-hw.mlir:20693:13
  wire            _T_424;	// matmul/matmul-hw.mlir:20676:13
  wire            _T_425;	// matmul/matmul-hw.mlir:20674:13
  wire            _T_426;	// matmul/matmul-hw.mlir:20673:13
  wire [31:0]     _T_427;	// matmul/matmul-hw.mlir:20664:13
  wire            _T_428;	// matmul/matmul-hw.mlir:20663:13
  wire            _T_429;	// matmul/matmul-hw.mlir:20646:13
  wire            _T_430;	// matmul/matmul-hw.mlir:20644:13
  wire            _T_431;	// matmul/matmul-hw.mlir:20643:13
  wire [31:0]     _T_432;	// matmul/matmul-hw.mlir:20642:13
  wire            _T_433;	// matmul/matmul-hw.mlir:20641:13
  wire [31:0]     _T_434;	// matmul/matmul-hw.mlir:20547:13
  wire            _T_435;	// matmul/matmul-hw.mlir:20546:13
  wire [3:0]      _T_436;	// matmul/matmul-hw.mlir:20545:13
  wire            _T_437;	// matmul/matmul-hw.mlir:20544:13
  wire            _T_438;	// matmul/matmul-hw.mlir:20528:13
  wire [31:0]     _T_439;	// matmul/matmul-hw.mlir:20519:13
  wire            _T_440;	// matmul/matmul-hw.mlir:20518:13
  wire            _T_441;	// matmul/matmul-hw.mlir:20501:13
  wire            _T_442;	// matmul/matmul-hw.mlir:20499:13
  wire            _T_443;	// matmul/matmul-hw.mlir:20498:13
  wire [31:0]     _T_444;	// matmul/matmul-hw.mlir:20489:13
  wire            _T_445;	// matmul/matmul-hw.mlir:20488:13
  wire            _T_446;	// matmul/matmul-hw.mlir:20471:13
  wire            _T_447;	// matmul/matmul-hw.mlir:20469:13
  wire            _T_448;	// matmul/matmul-hw.mlir:20468:13
  wire [31:0]     _T_449;	// matmul/matmul-hw.mlir:20459:13
  wire            _T_450;	// matmul/matmul-hw.mlir:20458:13
  wire            _T_451;	// matmul/matmul-hw.mlir:20441:13
  wire            _T_452;	// matmul/matmul-hw.mlir:20439:13
  wire            _T_453;	// matmul/matmul-hw.mlir:20438:13
  wire [31:0]     _T_454;	// matmul/matmul-hw.mlir:20429:13
  wire            _T_455;	// matmul/matmul-hw.mlir:20428:13
  wire            _T_456;	// matmul/matmul-hw.mlir:20411:13
  wire            _T_457;	// matmul/matmul-hw.mlir:20409:13
  wire            _T_458;	// matmul/matmul-hw.mlir:20408:13
  wire [31:0]     _T_459;	// matmul/matmul-hw.mlir:20399:13
  wire            _T_460;	// matmul/matmul-hw.mlir:20398:13
  wire            _T_461;	// matmul/matmul-hw.mlir:20381:13
  wire            _T_462;	// matmul/matmul-hw.mlir:20379:13
  wire            _T_463;	// matmul/matmul-hw.mlir:20378:13
  wire [31:0]     _T_464;	// matmul/matmul-hw.mlir:20369:13
  wire            _T_465;	// matmul/matmul-hw.mlir:20368:13
  wire            _T_466;	// matmul/matmul-hw.mlir:20351:13
  wire            _T_467;	// matmul/matmul-hw.mlir:20349:13
  wire            _T_468;	// matmul/matmul-hw.mlir:20348:13
  wire [31:0]     _T_469;	// matmul/matmul-hw.mlir:20339:13
  wire            _T_470;	// matmul/matmul-hw.mlir:20338:13
  wire            _T_471;	// matmul/matmul-hw.mlir:20321:13
  wire            _T_472;	// matmul/matmul-hw.mlir:20319:13
  wire            _T_473;	// matmul/matmul-hw.mlir:20318:13
  wire [31:0]     _T_474;	// matmul/matmul-hw.mlir:20309:13
  wire            _T_475;	// matmul/matmul-hw.mlir:20308:13
  wire            _T_476;	// matmul/matmul-hw.mlir:20291:13
  wire            _T_477;	// matmul/matmul-hw.mlir:20289:13
  wire            _T_478;	// matmul/matmul-hw.mlir:20288:13
  wire [31:0]     _T_479;	// matmul/matmul-hw.mlir:20279:13
  wire            _T_480;	// matmul/matmul-hw.mlir:20278:13
  wire            _T_481;	// matmul/matmul-hw.mlir:20261:13
  wire            _T_482;	// matmul/matmul-hw.mlir:20259:13
  wire            _T_483;	// matmul/matmul-hw.mlir:20258:13
  wire [31:0]     _T_484;	// matmul/matmul-hw.mlir:20249:13
  wire            _T_485;	// matmul/matmul-hw.mlir:20248:13
  wire            _T_486;	// matmul/matmul-hw.mlir:20231:13
  wire            _T_487;	// matmul/matmul-hw.mlir:20229:13
  wire            _T_488;	// matmul/matmul-hw.mlir:20228:13
  wire [31:0]     _T_489;	// matmul/matmul-hw.mlir:20219:13
  wire            _T_490;	// matmul/matmul-hw.mlir:20218:13
  wire            _T_491;	// matmul/matmul-hw.mlir:20201:13
  wire            _T_492;	// matmul/matmul-hw.mlir:20199:13
  wire            _T_493;	// matmul/matmul-hw.mlir:20198:13
  wire [31:0]     _T_494;	// matmul/matmul-hw.mlir:20189:13
  wire            _T_495;	// matmul/matmul-hw.mlir:20188:13
  wire            _T_496;	// matmul/matmul-hw.mlir:20171:13
  wire            _T_497;	// matmul/matmul-hw.mlir:20169:13
  wire            _T_498;	// matmul/matmul-hw.mlir:20168:13
  wire [31:0]     _T_499;	// matmul/matmul-hw.mlir:20159:13
  wire            _T_500;	// matmul/matmul-hw.mlir:20158:13
  wire            _T_501;	// matmul/matmul-hw.mlir:20141:13
  wire            _T_502;	// matmul/matmul-hw.mlir:20139:13
  wire            _T_503;	// matmul/matmul-hw.mlir:20138:13
  wire [31:0]     _T_504;	// matmul/matmul-hw.mlir:20129:13
  wire            _T_505;	// matmul/matmul-hw.mlir:20128:13
  wire            _T_506;	// matmul/matmul-hw.mlir:20111:13
  wire            _T_507;	// matmul/matmul-hw.mlir:20109:13
  wire            _T_508;	// matmul/matmul-hw.mlir:20108:13
  wire [31:0]     _T_509;	// matmul/matmul-hw.mlir:20099:13
  wire            _T_510;	// matmul/matmul-hw.mlir:20098:13
  wire            _T_511;	// matmul/matmul-hw.mlir:20081:13
  wire            _T_512;	// matmul/matmul-hw.mlir:20079:13
  wire            _T_513;	// matmul/matmul-hw.mlir:20078:13
  wire [31:0]     _T_514;	// matmul/matmul-hw.mlir:20069:13
  wire            _T_515;	// matmul/matmul-hw.mlir:20068:13
  wire            _T_516;	// matmul/matmul-hw.mlir:20051:13
  wire            _T_517;	// matmul/matmul-hw.mlir:20049:13
  wire            _T_518;	// matmul/matmul-hw.mlir:20048:13
  wire [31:0]     _T_519;	// matmul/matmul-hw.mlir:20047:13
  wire            _T_520;	// matmul/matmul-hw.mlir:20046:13
  wire [31:0]     _T_521;	// matmul/matmul-hw.mlir:19952:13
  wire            _T_522;	// matmul/matmul-hw.mlir:19951:13
  wire [3:0]      _T_523;	// matmul/matmul-hw.mlir:19950:13
  wire            _T_524;	// matmul/matmul-hw.mlir:19949:13
  wire            _T_525;	// matmul/matmul-hw.mlir:19933:13
  wire [31:0]     _T_526;	// matmul/matmul-hw.mlir:19924:13
  wire            _T_527;	// matmul/matmul-hw.mlir:19923:13
  wire            _T_528;	// matmul/matmul-hw.mlir:19906:13
  wire            _T_529;	// matmul/matmul-hw.mlir:19904:13
  wire            _T_530;	// matmul/matmul-hw.mlir:19903:13
  wire [31:0]     _T_531;	// matmul/matmul-hw.mlir:19894:13
  wire            _T_532;	// matmul/matmul-hw.mlir:19893:13
  wire            _T_533;	// matmul/matmul-hw.mlir:19876:13
  wire            _T_534;	// matmul/matmul-hw.mlir:19874:13
  wire            _T_535;	// matmul/matmul-hw.mlir:19873:13
  wire [31:0]     _T_536;	// matmul/matmul-hw.mlir:19864:13
  wire            _T_537;	// matmul/matmul-hw.mlir:19863:13
  wire            _T_538;	// matmul/matmul-hw.mlir:19846:13
  wire            _T_539;	// matmul/matmul-hw.mlir:19844:13
  wire            _T_540;	// matmul/matmul-hw.mlir:19843:13
  wire [31:0]     _T_541;	// matmul/matmul-hw.mlir:19834:13
  wire            _T_542;	// matmul/matmul-hw.mlir:19833:13
  wire            _T_543;	// matmul/matmul-hw.mlir:19816:13
  wire            _T_544;	// matmul/matmul-hw.mlir:19814:13
  wire            _T_545;	// matmul/matmul-hw.mlir:19813:13
  wire [31:0]     _T_546;	// matmul/matmul-hw.mlir:19804:13
  wire            _T_547;	// matmul/matmul-hw.mlir:19803:13
  wire            _T_548;	// matmul/matmul-hw.mlir:19786:13
  wire            _T_549;	// matmul/matmul-hw.mlir:19784:13
  wire            _T_550;	// matmul/matmul-hw.mlir:19783:13
  wire [31:0]     _T_551;	// matmul/matmul-hw.mlir:19774:13
  wire            _T_552;	// matmul/matmul-hw.mlir:19773:13
  wire            _T_553;	// matmul/matmul-hw.mlir:19756:13
  wire            _T_554;	// matmul/matmul-hw.mlir:19754:13
  wire            _T_555;	// matmul/matmul-hw.mlir:19753:13
  wire [31:0]     _T_556;	// matmul/matmul-hw.mlir:19744:13
  wire            _T_557;	// matmul/matmul-hw.mlir:19743:13
  wire            _T_558;	// matmul/matmul-hw.mlir:19726:13
  wire            _T_559;	// matmul/matmul-hw.mlir:19724:13
  wire            _T_560;	// matmul/matmul-hw.mlir:19723:13
  wire [31:0]     _T_561;	// matmul/matmul-hw.mlir:19714:13
  wire            _T_562;	// matmul/matmul-hw.mlir:19713:13
  wire            _T_563;	// matmul/matmul-hw.mlir:19696:13
  wire            _T_564;	// matmul/matmul-hw.mlir:19694:13
  wire            _T_565;	// matmul/matmul-hw.mlir:19693:13
  wire [31:0]     _T_566;	// matmul/matmul-hw.mlir:19684:13
  wire            _T_567;	// matmul/matmul-hw.mlir:19683:13
  wire            _T_568;	// matmul/matmul-hw.mlir:19666:13
  wire            _T_569;	// matmul/matmul-hw.mlir:19664:13
  wire            _T_570;	// matmul/matmul-hw.mlir:19663:13
  wire [31:0]     _T_571;	// matmul/matmul-hw.mlir:19654:13
  wire            _T_572;	// matmul/matmul-hw.mlir:19653:13
  wire            _T_573;	// matmul/matmul-hw.mlir:19636:13
  wire            _T_574;	// matmul/matmul-hw.mlir:19634:13
  wire            _T_575;	// matmul/matmul-hw.mlir:19633:13
  wire [31:0]     _T_576;	// matmul/matmul-hw.mlir:19624:13
  wire            _T_577;	// matmul/matmul-hw.mlir:19623:13
  wire            _T_578;	// matmul/matmul-hw.mlir:19606:13
  wire            _T_579;	// matmul/matmul-hw.mlir:19604:13
  wire            _T_580;	// matmul/matmul-hw.mlir:19603:13
  wire [31:0]     _T_581;	// matmul/matmul-hw.mlir:19594:13
  wire            _T_582;	// matmul/matmul-hw.mlir:19593:13
  wire            _T_583;	// matmul/matmul-hw.mlir:19576:13
  wire            _T_584;	// matmul/matmul-hw.mlir:19574:13
  wire            _T_585;	// matmul/matmul-hw.mlir:19573:13
  wire [31:0]     _T_586;	// matmul/matmul-hw.mlir:19564:13
  wire            _T_587;	// matmul/matmul-hw.mlir:19563:13
  wire            _T_588;	// matmul/matmul-hw.mlir:19546:13
  wire            _T_589;	// matmul/matmul-hw.mlir:19544:13
  wire            _T_590;	// matmul/matmul-hw.mlir:19543:13
  wire [31:0]     _T_591;	// matmul/matmul-hw.mlir:19534:13
  wire            _T_592;	// matmul/matmul-hw.mlir:19533:13
  wire            _T_593;	// matmul/matmul-hw.mlir:19516:13
  wire            _T_594;	// matmul/matmul-hw.mlir:19514:13
  wire            _T_595;	// matmul/matmul-hw.mlir:19513:13
  wire [31:0]     _T_596;	// matmul/matmul-hw.mlir:19504:13
  wire            _T_597;	// matmul/matmul-hw.mlir:19503:13
  wire            _T_598;	// matmul/matmul-hw.mlir:19486:13
  wire            _T_599;	// matmul/matmul-hw.mlir:19484:13
  wire            _T_600;	// matmul/matmul-hw.mlir:19483:13
  wire [31:0]     _T_601;	// matmul/matmul-hw.mlir:19474:13
  wire            _T_602;	// matmul/matmul-hw.mlir:19473:13
  wire            _T_603;	// matmul/matmul-hw.mlir:19456:13
  wire            _T_604;	// matmul/matmul-hw.mlir:19454:13
  wire            _T_605;	// matmul/matmul-hw.mlir:19453:13
  wire [31:0]     _T_606;	// matmul/matmul-hw.mlir:19452:13
  wire            _T_607;	// matmul/matmul-hw.mlir:19451:13
  wire [31:0]     _T_608;	// matmul/matmul-hw.mlir:19357:13
  wire            _T_609;	// matmul/matmul-hw.mlir:19356:13
  wire [3:0]      _T_610;	// matmul/matmul-hw.mlir:19355:13
  wire            _T_611;	// matmul/matmul-hw.mlir:19354:13
  wire            _T_612;	// matmul/matmul-hw.mlir:19338:13
  wire [31:0]     _T_613;	// matmul/matmul-hw.mlir:19329:13
  wire            _T_614;	// matmul/matmul-hw.mlir:19328:13
  wire            _T_615;	// matmul/matmul-hw.mlir:19311:13
  wire            _T_616;	// matmul/matmul-hw.mlir:19309:13
  wire            _T_617;	// matmul/matmul-hw.mlir:19308:13
  wire [31:0]     _T_618;	// matmul/matmul-hw.mlir:19299:13
  wire            _T_619;	// matmul/matmul-hw.mlir:19298:13
  wire            _T_620;	// matmul/matmul-hw.mlir:19281:13
  wire            _T_621;	// matmul/matmul-hw.mlir:19279:13
  wire            _T_622;	// matmul/matmul-hw.mlir:19278:13
  wire [31:0]     _T_623;	// matmul/matmul-hw.mlir:19269:13
  wire            _T_624;	// matmul/matmul-hw.mlir:19268:13
  wire            _T_625;	// matmul/matmul-hw.mlir:19251:13
  wire            _T_626;	// matmul/matmul-hw.mlir:19249:13
  wire            _T_627;	// matmul/matmul-hw.mlir:19248:13
  wire [31:0]     _T_628;	// matmul/matmul-hw.mlir:19239:13
  wire            _T_629;	// matmul/matmul-hw.mlir:19238:13
  wire            _T_630;	// matmul/matmul-hw.mlir:19221:13
  wire            _T_631;	// matmul/matmul-hw.mlir:19219:13
  wire            _T_632;	// matmul/matmul-hw.mlir:19218:13
  wire [31:0]     _T_633;	// matmul/matmul-hw.mlir:19209:13
  wire            _T_634;	// matmul/matmul-hw.mlir:19208:13
  wire            _T_635;	// matmul/matmul-hw.mlir:19191:13
  wire            _T_636;	// matmul/matmul-hw.mlir:19189:13
  wire            _T_637;	// matmul/matmul-hw.mlir:19188:13
  wire [31:0]     _T_638;	// matmul/matmul-hw.mlir:19179:13
  wire            _T_639;	// matmul/matmul-hw.mlir:19178:13
  wire            _T_640;	// matmul/matmul-hw.mlir:19161:13
  wire            _T_641;	// matmul/matmul-hw.mlir:19159:13
  wire            _T_642;	// matmul/matmul-hw.mlir:19158:13
  wire [31:0]     _T_643;	// matmul/matmul-hw.mlir:19149:13
  wire            _T_644;	// matmul/matmul-hw.mlir:19148:13
  wire            _T_645;	// matmul/matmul-hw.mlir:19131:13
  wire            _T_646;	// matmul/matmul-hw.mlir:19129:13
  wire            _T_647;	// matmul/matmul-hw.mlir:19128:13
  wire [31:0]     _T_648;	// matmul/matmul-hw.mlir:19119:13
  wire            _T_649;	// matmul/matmul-hw.mlir:19118:13
  wire            _T_650;	// matmul/matmul-hw.mlir:19101:13
  wire            _T_651;	// matmul/matmul-hw.mlir:19099:13
  wire            _T_652;	// matmul/matmul-hw.mlir:19098:13
  wire [31:0]     _T_653;	// matmul/matmul-hw.mlir:19089:13
  wire            _T_654;	// matmul/matmul-hw.mlir:19088:13
  wire            _T_655;	// matmul/matmul-hw.mlir:19071:13
  wire            _T_656;	// matmul/matmul-hw.mlir:19069:13
  wire            _T_657;	// matmul/matmul-hw.mlir:19068:13
  wire [31:0]     _T_658;	// matmul/matmul-hw.mlir:19059:13
  wire            _T_659;	// matmul/matmul-hw.mlir:19058:13
  wire            _T_660;	// matmul/matmul-hw.mlir:19041:13
  wire            _T_661;	// matmul/matmul-hw.mlir:19039:13
  wire            _T_662;	// matmul/matmul-hw.mlir:19038:13
  wire [31:0]     _T_663;	// matmul/matmul-hw.mlir:19029:13
  wire            _T_664;	// matmul/matmul-hw.mlir:19028:13
  wire            _T_665;	// matmul/matmul-hw.mlir:19011:13
  wire            _T_666;	// matmul/matmul-hw.mlir:19009:13
  wire            _T_667;	// matmul/matmul-hw.mlir:19008:13
  wire [31:0]     _T_668;	// matmul/matmul-hw.mlir:18999:13
  wire            _T_669;	// matmul/matmul-hw.mlir:18998:13
  wire            _T_670;	// matmul/matmul-hw.mlir:18981:13
  wire            _T_671;	// matmul/matmul-hw.mlir:18979:13
  wire            _T_672;	// matmul/matmul-hw.mlir:18978:13
  wire [31:0]     _T_673;	// matmul/matmul-hw.mlir:18969:13
  wire            _T_674;	// matmul/matmul-hw.mlir:18968:13
  wire            _T_675;	// matmul/matmul-hw.mlir:18951:13
  wire            _T_676;	// matmul/matmul-hw.mlir:18949:13
  wire            _T_677;	// matmul/matmul-hw.mlir:18948:13
  wire [31:0]     _T_678;	// matmul/matmul-hw.mlir:18939:13
  wire            _T_679;	// matmul/matmul-hw.mlir:18938:13
  wire            _T_680;	// matmul/matmul-hw.mlir:18921:13
  wire            _T_681;	// matmul/matmul-hw.mlir:18919:13
  wire            _T_682;	// matmul/matmul-hw.mlir:18918:13
  wire [31:0]     _T_683;	// matmul/matmul-hw.mlir:18909:13
  wire            _T_684;	// matmul/matmul-hw.mlir:18908:13
  wire            _T_685;	// matmul/matmul-hw.mlir:18891:13
  wire            _T_686;	// matmul/matmul-hw.mlir:18889:13
  wire            _T_687;	// matmul/matmul-hw.mlir:18888:13
  wire [31:0]     _T_688;	// matmul/matmul-hw.mlir:18879:13
  wire            _T_689;	// matmul/matmul-hw.mlir:18878:13
  wire            _T_690;	// matmul/matmul-hw.mlir:18861:13
  wire            _T_691;	// matmul/matmul-hw.mlir:18859:13
  wire            _T_692;	// matmul/matmul-hw.mlir:18858:13
  wire [31:0]     _T_693;	// matmul/matmul-hw.mlir:18857:13
  wire            _T_694;	// matmul/matmul-hw.mlir:18856:13
  wire [31:0]     _T_695;	// matmul/matmul-hw.mlir:18762:13
  wire            _T_696;	// matmul/matmul-hw.mlir:18761:13
  wire [3:0]      _T_697;	// matmul/matmul-hw.mlir:18760:13
  wire            _T_698;	// matmul/matmul-hw.mlir:18759:13
  wire            _T_699;	// matmul/matmul-hw.mlir:18743:13
  wire [31:0]     _T_700;	// matmul/matmul-hw.mlir:18734:13
  wire            _T_701;	// matmul/matmul-hw.mlir:18733:13
  wire            _T_702;	// matmul/matmul-hw.mlir:18716:13
  wire            _T_703;	// matmul/matmul-hw.mlir:18714:13
  wire            _T_704;	// matmul/matmul-hw.mlir:18713:13
  wire [31:0]     _T_705;	// matmul/matmul-hw.mlir:18704:13
  wire            _T_706;	// matmul/matmul-hw.mlir:18703:13
  wire            _T_707;	// matmul/matmul-hw.mlir:18686:13
  wire            _T_708;	// matmul/matmul-hw.mlir:18684:13
  wire            _T_709;	// matmul/matmul-hw.mlir:18683:13
  wire [31:0]     _T_710;	// matmul/matmul-hw.mlir:18674:13
  wire            _T_711;	// matmul/matmul-hw.mlir:18673:13
  wire            _T_712;	// matmul/matmul-hw.mlir:18656:13
  wire            _T_713;	// matmul/matmul-hw.mlir:18654:13
  wire            _T_714;	// matmul/matmul-hw.mlir:18653:13
  wire [31:0]     _T_715;	// matmul/matmul-hw.mlir:18644:13
  wire            _T_716;	// matmul/matmul-hw.mlir:18643:13
  wire            _T_717;	// matmul/matmul-hw.mlir:18626:13
  wire            _T_718;	// matmul/matmul-hw.mlir:18624:13
  wire            _T_719;	// matmul/matmul-hw.mlir:18623:13
  wire [31:0]     _T_720;	// matmul/matmul-hw.mlir:18614:13
  wire            _T_721;	// matmul/matmul-hw.mlir:18613:13
  wire            _T_722;	// matmul/matmul-hw.mlir:18596:13
  wire            _T_723;	// matmul/matmul-hw.mlir:18594:13
  wire            _T_724;	// matmul/matmul-hw.mlir:18593:13
  wire [31:0]     _T_725;	// matmul/matmul-hw.mlir:18584:13
  wire            _T_726;	// matmul/matmul-hw.mlir:18583:13
  wire            _T_727;	// matmul/matmul-hw.mlir:18566:13
  wire            _T_728;	// matmul/matmul-hw.mlir:18564:13
  wire            _T_729;	// matmul/matmul-hw.mlir:18563:13
  wire [31:0]     _T_730;	// matmul/matmul-hw.mlir:18554:13
  wire            _T_731;	// matmul/matmul-hw.mlir:18553:13
  wire            _T_732;	// matmul/matmul-hw.mlir:18536:13
  wire            _T_733;	// matmul/matmul-hw.mlir:18534:13
  wire            _T_734;	// matmul/matmul-hw.mlir:18533:13
  wire [31:0]     _T_735;	// matmul/matmul-hw.mlir:18524:13
  wire            _T_736;	// matmul/matmul-hw.mlir:18523:13
  wire            _T_737;	// matmul/matmul-hw.mlir:18506:13
  wire            _T_738;	// matmul/matmul-hw.mlir:18504:13
  wire            _T_739;	// matmul/matmul-hw.mlir:18503:13
  wire [31:0]     _T_740;	// matmul/matmul-hw.mlir:18494:13
  wire            _T_741;	// matmul/matmul-hw.mlir:18493:13
  wire            _T_742;	// matmul/matmul-hw.mlir:18476:13
  wire            _T_743;	// matmul/matmul-hw.mlir:18474:13
  wire            _T_744;	// matmul/matmul-hw.mlir:18473:13
  wire [31:0]     _T_745;	// matmul/matmul-hw.mlir:18464:13
  wire            _T_746;	// matmul/matmul-hw.mlir:18463:13
  wire            _T_747;	// matmul/matmul-hw.mlir:18446:13
  wire            _T_748;	// matmul/matmul-hw.mlir:18444:13
  wire            _T_749;	// matmul/matmul-hw.mlir:18443:13
  wire [31:0]     _T_750;	// matmul/matmul-hw.mlir:18434:13
  wire            _T_751;	// matmul/matmul-hw.mlir:18433:13
  wire            _T_752;	// matmul/matmul-hw.mlir:18416:13
  wire            _T_753;	// matmul/matmul-hw.mlir:18414:13
  wire            _T_754;	// matmul/matmul-hw.mlir:18413:13
  wire [31:0]     _T_755;	// matmul/matmul-hw.mlir:18404:13
  wire            _T_756;	// matmul/matmul-hw.mlir:18403:13
  wire            _T_757;	// matmul/matmul-hw.mlir:18386:13
  wire            _T_758;	// matmul/matmul-hw.mlir:18384:13
  wire            _T_759;	// matmul/matmul-hw.mlir:18383:13
  wire [31:0]     _T_760;	// matmul/matmul-hw.mlir:18374:13
  wire            _T_761;	// matmul/matmul-hw.mlir:18373:13
  wire            _T_762;	// matmul/matmul-hw.mlir:18356:13
  wire            _T_763;	// matmul/matmul-hw.mlir:18354:13
  wire            _T_764;	// matmul/matmul-hw.mlir:18353:13
  wire [31:0]     _T_765;	// matmul/matmul-hw.mlir:18344:13
  wire            _T_766;	// matmul/matmul-hw.mlir:18343:13
  wire            _T_767;	// matmul/matmul-hw.mlir:18326:13
  wire            _T_768;	// matmul/matmul-hw.mlir:18324:13
  wire            _T_769;	// matmul/matmul-hw.mlir:18323:13
  wire [31:0]     _T_770;	// matmul/matmul-hw.mlir:18314:13
  wire            _T_771;	// matmul/matmul-hw.mlir:18313:13
  wire            _T_772;	// matmul/matmul-hw.mlir:18296:13
  wire            _T_773;	// matmul/matmul-hw.mlir:18294:13
  wire            _T_774;	// matmul/matmul-hw.mlir:18293:13
  wire [31:0]     _T_775;	// matmul/matmul-hw.mlir:18284:13
  wire            _T_776;	// matmul/matmul-hw.mlir:18283:13
  wire            _T_777;	// matmul/matmul-hw.mlir:18266:13
  wire            _T_778;	// matmul/matmul-hw.mlir:18264:13
  wire            _T_779;	// matmul/matmul-hw.mlir:18263:13
  wire [31:0]     _T_780;	// matmul/matmul-hw.mlir:18262:13
  wire            _T_781;	// matmul/matmul-hw.mlir:18261:13
  wire [31:0]     _T_782;	// matmul/matmul-hw.mlir:18167:13
  wire            _T_783;	// matmul/matmul-hw.mlir:18166:13
  wire [3:0]      _T_784;	// matmul/matmul-hw.mlir:18165:13
  wire            _T_785;	// matmul/matmul-hw.mlir:18164:13
  wire            _T_786;	// matmul/matmul-hw.mlir:18148:13
  wire [31:0]     _T_787;	// matmul/matmul-hw.mlir:18139:13
  wire            _T_788;	// matmul/matmul-hw.mlir:18138:13
  wire            _T_789;	// matmul/matmul-hw.mlir:18121:13
  wire            _T_790;	// matmul/matmul-hw.mlir:18119:13
  wire            _T_791;	// matmul/matmul-hw.mlir:18118:13
  wire [31:0]     _T_792;	// matmul/matmul-hw.mlir:18109:13
  wire            _T_793;	// matmul/matmul-hw.mlir:18108:13
  wire            _T_794;	// matmul/matmul-hw.mlir:18091:13
  wire            _T_795;	// matmul/matmul-hw.mlir:18089:13
  wire            _T_796;	// matmul/matmul-hw.mlir:18088:13
  wire [31:0]     _T_797;	// matmul/matmul-hw.mlir:18079:13
  wire            _T_798;	// matmul/matmul-hw.mlir:18078:13
  wire            _T_799;	// matmul/matmul-hw.mlir:18061:13
  wire            _T_800;	// matmul/matmul-hw.mlir:18059:13
  wire            _T_801;	// matmul/matmul-hw.mlir:18058:13
  wire [31:0]     _T_802;	// matmul/matmul-hw.mlir:18049:13
  wire            _T_803;	// matmul/matmul-hw.mlir:18048:13
  wire            _T_804;	// matmul/matmul-hw.mlir:18031:13
  wire            _T_805;	// matmul/matmul-hw.mlir:18029:13
  wire            _T_806;	// matmul/matmul-hw.mlir:18028:13
  wire [31:0]     _T_807;	// matmul/matmul-hw.mlir:18019:13
  wire            _T_808;	// matmul/matmul-hw.mlir:18018:13
  wire            _T_809;	// matmul/matmul-hw.mlir:18001:13
  wire            _T_810;	// matmul/matmul-hw.mlir:17999:13
  wire            _T_811;	// matmul/matmul-hw.mlir:17998:13
  wire [31:0]     _T_812;	// matmul/matmul-hw.mlir:17989:13
  wire            _T_813;	// matmul/matmul-hw.mlir:17988:13
  wire            _T_814;	// matmul/matmul-hw.mlir:17971:13
  wire            _T_815;	// matmul/matmul-hw.mlir:17969:13
  wire            _T_816;	// matmul/matmul-hw.mlir:17968:13
  wire [31:0]     _T_817;	// matmul/matmul-hw.mlir:17959:13
  wire            _T_818;	// matmul/matmul-hw.mlir:17958:13
  wire            _T_819;	// matmul/matmul-hw.mlir:17941:13
  wire            _T_820;	// matmul/matmul-hw.mlir:17939:13
  wire            _T_821;	// matmul/matmul-hw.mlir:17938:13
  wire [31:0]     _T_822;	// matmul/matmul-hw.mlir:17929:13
  wire            _T_823;	// matmul/matmul-hw.mlir:17928:13
  wire            _T_824;	// matmul/matmul-hw.mlir:17911:13
  wire            _T_825;	// matmul/matmul-hw.mlir:17909:13
  wire            _T_826;	// matmul/matmul-hw.mlir:17908:13
  wire [31:0]     _T_827;	// matmul/matmul-hw.mlir:17899:13
  wire            _T_828;	// matmul/matmul-hw.mlir:17898:13
  wire            _T_829;	// matmul/matmul-hw.mlir:17881:13
  wire            _T_830;	// matmul/matmul-hw.mlir:17879:13
  wire            _T_831;	// matmul/matmul-hw.mlir:17878:13
  wire [31:0]     _T_832;	// matmul/matmul-hw.mlir:17869:13
  wire            _T_833;	// matmul/matmul-hw.mlir:17868:13
  wire            _T_834;	// matmul/matmul-hw.mlir:17851:13
  wire            _T_835;	// matmul/matmul-hw.mlir:17849:13
  wire            _T_836;	// matmul/matmul-hw.mlir:17848:13
  wire [31:0]     _T_837;	// matmul/matmul-hw.mlir:17839:13
  wire            _T_838;	// matmul/matmul-hw.mlir:17838:13
  wire            _T_839;	// matmul/matmul-hw.mlir:17821:13
  wire            _T_840;	// matmul/matmul-hw.mlir:17819:13
  wire            _T_841;	// matmul/matmul-hw.mlir:17818:13
  wire [31:0]     _T_842;	// matmul/matmul-hw.mlir:17809:13
  wire            _T_843;	// matmul/matmul-hw.mlir:17808:13
  wire            _T_844;	// matmul/matmul-hw.mlir:17791:13
  wire            _T_845;	// matmul/matmul-hw.mlir:17789:13
  wire            _T_846;	// matmul/matmul-hw.mlir:17788:13
  wire [31:0]     _T_847;	// matmul/matmul-hw.mlir:17779:13
  wire            _T_848;	// matmul/matmul-hw.mlir:17778:13
  wire            _T_849;	// matmul/matmul-hw.mlir:17761:13
  wire            _T_850;	// matmul/matmul-hw.mlir:17759:13
  wire            _T_851;	// matmul/matmul-hw.mlir:17758:13
  wire [31:0]     _T_852;	// matmul/matmul-hw.mlir:17749:13
  wire            _T_853;	// matmul/matmul-hw.mlir:17748:13
  wire            _T_854;	// matmul/matmul-hw.mlir:17731:13
  wire            _T_855;	// matmul/matmul-hw.mlir:17729:13
  wire            _T_856;	// matmul/matmul-hw.mlir:17728:13
  wire [31:0]     _T_857;	// matmul/matmul-hw.mlir:17719:13
  wire            _T_858;	// matmul/matmul-hw.mlir:17718:13
  wire            _T_859;	// matmul/matmul-hw.mlir:17701:13
  wire            _T_860;	// matmul/matmul-hw.mlir:17699:13
  wire            _T_861;	// matmul/matmul-hw.mlir:17698:13
  wire [31:0]     _T_862;	// matmul/matmul-hw.mlir:17689:13
  wire            _T_863;	// matmul/matmul-hw.mlir:17688:13
  wire            _T_864;	// matmul/matmul-hw.mlir:17671:13
  wire            _T_865;	// matmul/matmul-hw.mlir:17669:13
  wire            _T_866;	// matmul/matmul-hw.mlir:17668:13
  wire [31:0]     _T_867;	// matmul/matmul-hw.mlir:17667:13
  wire            _T_868;	// matmul/matmul-hw.mlir:17666:13
  wire [31:0]     _T_869;	// matmul/matmul-hw.mlir:17572:13
  wire            _T_870;	// matmul/matmul-hw.mlir:17571:13
  wire [3:0]      _T_871;	// matmul/matmul-hw.mlir:17570:13
  wire            _T_872;	// matmul/matmul-hw.mlir:17569:13
  wire            _T_873;	// matmul/matmul-hw.mlir:17553:13
  wire [31:0]     _T_874;	// matmul/matmul-hw.mlir:17544:13
  wire            _T_875;	// matmul/matmul-hw.mlir:17543:13
  wire            _T_876;	// matmul/matmul-hw.mlir:17526:13
  wire            _T_877;	// matmul/matmul-hw.mlir:17524:13
  wire            _T_878;	// matmul/matmul-hw.mlir:17523:13
  wire [31:0]     _T_879;	// matmul/matmul-hw.mlir:17514:13
  wire            _T_880;	// matmul/matmul-hw.mlir:17513:13
  wire            _T_881;	// matmul/matmul-hw.mlir:17496:13
  wire            _T_882;	// matmul/matmul-hw.mlir:17494:13
  wire            _T_883;	// matmul/matmul-hw.mlir:17493:13
  wire [31:0]     _T_884;	// matmul/matmul-hw.mlir:17484:13
  wire            _T_885;	// matmul/matmul-hw.mlir:17483:13
  wire            _T_886;	// matmul/matmul-hw.mlir:17466:13
  wire            _T_887;	// matmul/matmul-hw.mlir:17464:13
  wire            _T_888;	// matmul/matmul-hw.mlir:17463:13
  wire [31:0]     _T_889;	// matmul/matmul-hw.mlir:17454:13
  wire            _T_890;	// matmul/matmul-hw.mlir:17453:13
  wire            _T_891;	// matmul/matmul-hw.mlir:17436:13
  wire            _T_892;	// matmul/matmul-hw.mlir:17434:13
  wire            _T_893;	// matmul/matmul-hw.mlir:17433:13
  wire [31:0]     _T_894;	// matmul/matmul-hw.mlir:17424:13
  wire            _T_895;	// matmul/matmul-hw.mlir:17423:13
  wire            _T_896;	// matmul/matmul-hw.mlir:17406:13
  wire            _T_897;	// matmul/matmul-hw.mlir:17404:13
  wire            _T_898;	// matmul/matmul-hw.mlir:17403:13
  wire [31:0]     _T_899;	// matmul/matmul-hw.mlir:17394:13
  wire            _T_900;	// matmul/matmul-hw.mlir:17393:13
  wire            _T_901;	// matmul/matmul-hw.mlir:17376:13
  wire            _T_902;	// matmul/matmul-hw.mlir:17374:13
  wire            _T_903;	// matmul/matmul-hw.mlir:17373:13
  wire [31:0]     _T_904;	// matmul/matmul-hw.mlir:17364:13
  wire            _T_905;	// matmul/matmul-hw.mlir:17363:13
  wire            _T_906;	// matmul/matmul-hw.mlir:17346:13
  wire            _T_907;	// matmul/matmul-hw.mlir:17344:13
  wire            _T_908;	// matmul/matmul-hw.mlir:17343:13
  wire [31:0]     _T_909;	// matmul/matmul-hw.mlir:17334:13
  wire            _T_910;	// matmul/matmul-hw.mlir:17333:13
  wire            _T_911;	// matmul/matmul-hw.mlir:17316:13
  wire            _T_912;	// matmul/matmul-hw.mlir:17314:13
  wire            _T_913;	// matmul/matmul-hw.mlir:17313:13
  wire [31:0]     _T_914;	// matmul/matmul-hw.mlir:17304:13
  wire            _T_915;	// matmul/matmul-hw.mlir:17303:13
  wire            _T_916;	// matmul/matmul-hw.mlir:17286:13
  wire            _T_917;	// matmul/matmul-hw.mlir:17284:13
  wire            _T_918;	// matmul/matmul-hw.mlir:17283:13
  wire [31:0]     _T_919;	// matmul/matmul-hw.mlir:17274:13
  wire            _T_920;	// matmul/matmul-hw.mlir:17273:13
  wire            _T_921;	// matmul/matmul-hw.mlir:17256:13
  wire            _T_922;	// matmul/matmul-hw.mlir:17254:13
  wire            _T_923;	// matmul/matmul-hw.mlir:17253:13
  wire [31:0]     _T_924;	// matmul/matmul-hw.mlir:17244:13
  wire            _T_925;	// matmul/matmul-hw.mlir:17243:13
  wire            _T_926;	// matmul/matmul-hw.mlir:17226:13
  wire            _T_927;	// matmul/matmul-hw.mlir:17224:13
  wire            _T_928;	// matmul/matmul-hw.mlir:17223:13
  wire [31:0]     _T_929;	// matmul/matmul-hw.mlir:17214:13
  wire            _T_930;	// matmul/matmul-hw.mlir:17213:13
  wire            _T_931;	// matmul/matmul-hw.mlir:17196:13
  wire            _T_932;	// matmul/matmul-hw.mlir:17194:13
  wire            _T_933;	// matmul/matmul-hw.mlir:17193:13
  wire [31:0]     _T_934;	// matmul/matmul-hw.mlir:17184:13
  wire            _T_935;	// matmul/matmul-hw.mlir:17183:13
  wire            _T_936;	// matmul/matmul-hw.mlir:17166:13
  wire            _T_937;	// matmul/matmul-hw.mlir:17164:13
  wire            _T_938;	// matmul/matmul-hw.mlir:17163:13
  wire [31:0]     _T_939;	// matmul/matmul-hw.mlir:17154:13
  wire            _T_940;	// matmul/matmul-hw.mlir:17153:13
  wire            _T_941;	// matmul/matmul-hw.mlir:17136:13
  wire            _T_942;	// matmul/matmul-hw.mlir:17134:13
  wire            _T_943;	// matmul/matmul-hw.mlir:17133:13
  wire [31:0]     _T_944;	// matmul/matmul-hw.mlir:17124:13
  wire            _T_945;	// matmul/matmul-hw.mlir:17123:13
  wire            _T_946;	// matmul/matmul-hw.mlir:17106:13
  wire            _T_947;	// matmul/matmul-hw.mlir:17104:13
  wire            _T_948;	// matmul/matmul-hw.mlir:17103:13
  wire [31:0]     _T_949;	// matmul/matmul-hw.mlir:17094:13
  wire            _T_950;	// matmul/matmul-hw.mlir:17093:13
  wire            _T_951;	// matmul/matmul-hw.mlir:17076:13
  wire            _T_952;	// matmul/matmul-hw.mlir:17074:13
  wire            _T_953;	// matmul/matmul-hw.mlir:17073:13
  wire [31:0]     _T_954;	// matmul/matmul-hw.mlir:17072:13
  wire            _T_955;	// matmul/matmul-hw.mlir:17071:13
  wire [31:0]     _T_956;	// matmul/matmul-hw.mlir:16977:13
  wire            _T_957;	// matmul/matmul-hw.mlir:16976:13
  wire [3:0]      _T_958;	// matmul/matmul-hw.mlir:16975:13
  wire            _T_959;	// matmul/matmul-hw.mlir:16974:13
  wire            _T_960;	// matmul/matmul-hw.mlir:16958:13
  wire [31:0]     _T_961;	// matmul/matmul-hw.mlir:16949:13
  wire            _T_962;	// matmul/matmul-hw.mlir:16948:13
  wire            _T_963;	// matmul/matmul-hw.mlir:16931:13
  wire            _T_964;	// matmul/matmul-hw.mlir:16929:13
  wire            _T_965;	// matmul/matmul-hw.mlir:16928:13
  wire [31:0]     _T_966;	// matmul/matmul-hw.mlir:16919:13
  wire            _T_967;	// matmul/matmul-hw.mlir:16918:13
  wire            _T_968;	// matmul/matmul-hw.mlir:16901:13
  wire            _T_969;	// matmul/matmul-hw.mlir:16899:13
  wire            _T_970;	// matmul/matmul-hw.mlir:16898:13
  wire [31:0]     _T_971;	// matmul/matmul-hw.mlir:16889:13
  wire            _T_972;	// matmul/matmul-hw.mlir:16888:13
  wire            _T_973;	// matmul/matmul-hw.mlir:16871:13
  wire            _T_974;	// matmul/matmul-hw.mlir:16869:13
  wire            _T_975;	// matmul/matmul-hw.mlir:16868:13
  wire [31:0]     _T_976;	// matmul/matmul-hw.mlir:16859:13
  wire            _T_977;	// matmul/matmul-hw.mlir:16858:13
  wire            _T_978;	// matmul/matmul-hw.mlir:16841:13
  wire            _T_979;	// matmul/matmul-hw.mlir:16839:13
  wire            _T_980;	// matmul/matmul-hw.mlir:16838:13
  wire [31:0]     _T_981;	// matmul/matmul-hw.mlir:16829:13
  wire            _T_982;	// matmul/matmul-hw.mlir:16828:13
  wire            _T_983;	// matmul/matmul-hw.mlir:16811:13
  wire            _T_984;	// matmul/matmul-hw.mlir:16809:13
  wire            _T_985;	// matmul/matmul-hw.mlir:16808:13
  wire [31:0]     _T_986;	// matmul/matmul-hw.mlir:16799:13
  wire            _T_987;	// matmul/matmul-hw.mlir:16798:13
  wire            _T_988;	// matmul/matmul-hw.mlir:16781:13
  wire            _T_989;	// matmul/matmul-hw.mlir:16779:13
  wire            _T_990;	// matmul/matmul-hw.mlir:16778:13
  wire [31:0]     _T_991;	// matmul/matmul-hw.mlir:16769:13
  wire            _T_992;	// matmul/matmul-hw.mlir:16768:13
  wire            _T_993;	// matmul/matmul-hw.mlir:16751:13
  wire            _T_994;	// matmul/matmul-hw.mlir:16749:13
  wire            _T_995;	// matmul/matmul-hw.mlir:16748:13
  wire [31:0]     _T_996;	// matmul/matmul-hw.mlir:16739:13
  wire            _T_997;	// matmul/matmul-hw.mlir:16738:13
  wire            _T_998;	// matmul/matmul-hw.mlir:16721:13
  wire            _T_999;	// matmul/matmul-hw.mlir:16719:13
  wire            _T_1000;	// matmul/matmul-hw.mlir:16718:13
  wire [31:0]     _T_1001;	// matmul/matmul-hw.mlir:16709:13
  wire            _T_1002;	// matmul/matmul-hw.mlir:16708:13
  wire            _T_1003;	// matmul/matmul-hw.mlir:16691:13
  wire            _T_1004;	// matmul/matmul-hw.mlir:16689:13
  wire            _T_1005;	// matmul/matmul-hw.mlir:16688:13
  wire [31:0]     _T_1006;	// matmul/matmul-hw.mlir:16679:13
  wire            _T_1007;	// matmul/matmul-hw.mlir:16678:13
  wire            _T_1008;	// matmul/matmul-hw.mlir:16661:13
  wire            _T_1009;	// matmul/matmul-hw.mlir:16659:13
  wire            _T_1010;	// matmul/matmul-hw.mlir:16658:13
  wire [31:0]     _T_1011;	// matmul/matmul-hw.mlir:16649:13
  wire            _T_1012;	// matmul/matmul-hw.mlir:16648:13
  wire            _T_1013;	// matmul/matmul-hw.mlir:16631:13
  wire            _T_1014;	// matmul/matmul-hw.mlir:16629:13
  wire            _T_1015;	// matmul/matmul-hw.mlir:16628:13
  wire [31:0]     _T_1016;	// matmul/matmul-hw.mlir:16619:13
  wire            _T_1017;	// matmul/matmul-hw.mlir:16618:13
  wire            _T_1018;	// matmul/matmul-hw.mlir:16601:13
  wire            _T_1019;	// matmul/matmul-hw.mlir:16599:13
  wire            _T_1020;	// matmul/matmul-hw.mlir:16598:13
  wire [31:0]     _T_1021;	// matmul/matmul-hw.mlir:16589:13
  wire            _T_1022;	// matmul/matmul-hw.mlir:16588:13
  wire            _T_1023;	// matmul/matmul-hw.mlir:16571:13
  wire            _T_1024;	// matmul/matmul-hw.mlir:16569:13
  wire            _T_1025;	// matmul/matmul-hw.mlir:16568:13
  wire [31:0]     _T_1026;	// matmul/matmul-hw.mlir:16559:13
  wire            _T_1027;	// matmul/matmul-hw.mlir:16558:13
  wire            _T_1028;	// matmul/matmul-hw.mlir:16541:13
  wire            _T_1029;	// matmul/matmul-hw.mlir:16539:13
  wire            _T_1030;	// matmul/matmul-hw.mlir:16538:13
  wire [31:0]     _T_1031;	// matmul/matmul-hw.mlir:16529:13
  wire            _T_1032;	// matmul/matmul-hw.mlir:16528:13
  wire            _T_1033;	// matmul/matmul-hw.mlir:16511:13
  wire            _T_1034;	// matmul/matmul-hw.mlir:16509:13
  wire            _T_1035;	// matmul/matmul-hw.mlir:16508:13
  wire [31:0]     _T_1036;	// matmul/matmul-hw.mlir:16499:13
  wire            _T_1037;	// matmul/matmul-hw.mlir:16498:13
  wire            _T_1038;	// matmul/matmul-hw.mlir:16481:13
  wire            _T_1039;	// matmul/matmul-hw.mlir:16479:13
  wire            _T_1040;	// matmul/matmul-hw.mlir:16478:13
  wire [31:0]     _T_1041;	// matmul/matmul-hw.mlir:16477:13
  wire            _T_1042;	// matmul/matmul-hw.mlir:16476:13
  wire [31:0]     _T_1043;	// matmul/matmul-hw.mlir:16382:13
  wire            _T_1044;	// matmul/matmul-hw.mlir:16381:13
  wire [3:0]      _T_1045;	// matmul/matmul-hw.mlir:16380:13
  wire            _T_1046;	// matmul/matmul-hw.mlir:16379:13
  wire            _T_1047;	// matmul/matmul-hw.mlir:16363:13
  wire [31:0]     _T_1048;	// matmul/matmul-hw.mlir:16354:13
  wire            _T_1049;	// matmul/matmul-hw.mlir:16353:13
  wire            _T_1050;	// matmul/matmul-hw.mlir:16336:13
  wire            _T_1051;	// matmul/matmul-hw.mlir:16334:13
  wire            _T_1052;	// matmul/matmul-hw.mlir:16333:13
  wire [31:0]     _T_1053;	// matmul/matmul-hw.mlir:16324:13
  wire            _T_1054;	// matmul/matmul-hw.mlir:16323:13
  wire            _T_1055;	// matmul/matmul-hw.mlir:16306:13
  wire            _T_1056;	// matmul/matmul-hw.mlir:16304:13
  wire            _T_1057;	// matmul/matmul-hw.mlir:16303:13
  wire [31:0]     _T_1058;	// matmul/matmul-hw.mlir:16294:13
  wire            _T_1059;	// matmul/matmul-hw.mlir:16293:13
  wire            _T_1060;	// matmul/matmul-hw.mlir:16276:13
  wire            _T_1061;	// matmul/matmul-hw.mlir:16274:13
  wire            _T_1062;	// matmul/matmul-hw.mlir:16273:13
  wire [31:0]     _T_1063;	// matmul/matmul-hw.mlir:16264:13
  wire            _T_1064;	// matmul/matmul-hw.mlir:16263:13
  wire            _T_1065;	// matmul/matmul-hw.mlir:16246:13
  wire            _T_1066;	// matmul/matmul-hw.mlir:16244:13
  wire            _T_1067;	// matmul/matmul-hw.mlir:16243:13
  wire [31:0]     _T_1068;	// matmul/matmul-hw.mlir:16234:13
  wire            _T_1069;	// matmul/matmul-hw.mlir:16233:13
  wire            _T_1070;	// matmul/matmul-hw.mlir:16216:13
  wire            _T_1071;	// matmul/matmul-hw.mlir:16214:13
  wire            _T_1072;	// matmul/matmul-hw.mlir:16213:13
  wire [31:0]     _T_1073;	// matmul/matmul-hw.mlir:16204:13
  wire            _T_1074;	// matmul/matmul-hw.mlir:16203:13
  wire            _T_1075;	// matmul/matmul-hw.mlir:16186:13
  wire            _T_1076;	// matmul/matmul-hw.mlir:16184:13
  wire            _T_1077;	// matmul/matmul-hw.mlir:16183:13
  wire [31:0]     _T_1078;	// matmul/matmul-hw.mlir:16174:13
  wire            _T_1079;	// matmul/matmul-hw.mlir:16173:13
  wire            _T_1080;	// matmul/matmul-hw.mlir:16156:13
  wire            _T_1081;	// matmul/matmul-hw.mlir:16154:13
  wire            _T_1082;	// matmul/matmul-hw.mlir:16153:13
  wire [31:0]     _T_1083;	// matmul/matmul-hw.mlir:16144:13
  wire            _T_1084;	// matmul/matmul-hw.mlir:16143:13
  wire            _T_1085;	// matmul/matmul-hw.mlir:16126:13
  wire            _T_1086;	// matmul/matmul-hw.mlir:16124:13
  wire            _T_1087;	// matmul/matmul-hw.mlir:16123:13
  wire [31:0]     _T_1088;	// matmul/matmul-hw.mlir:16114:13
  wire            _T_1089;	// matmul/matmul-hw.mlir:16113:13
  wire            _T_1090;	// matmul/matmul-hw.mlir:16096:13
  wire            _T_1091;	// matmul/matmul-hw.mlir:16094:13
  wire            _T_1092;	// matmul/matmul-hw.mlir:16093:13
  wire [31:0]     _T_1093;	// matmul/matmul-hw.mlir:16084:13
  wire            _T_1094;	// matmul/matmul-hw.mlir:16083:13
  wire            _T_1095;	// matmul/matmul-hw.mlir:16066:13
  wire            _T_1096;	// matmul/matmul-hw.mlir:16064:13
  wire            _T_1097;	// matmul/matmul-hw.mlir:16063:13
  wire [31:0]     _T_1098;	// matmul/matmul-hw.mlir:16054:13
  wire            _T_1099;	// matmul/matmul-hw.mlir:16053:13
  wire            _T_1100;	// matmul/matmul-hw.mlir:16036:13
  wire            _T_1101;	// matmul/matmul-hw.mlir:16034:13
  wire            _T_1102;	// matmul/matmul-hw.mlir:16033:13
  wire [31:0]     _T_1103;	// matmul/matmul-hw.mlir:16024:13
  wire            _T_1104;	// matmul/matmul-hw.mlir:16023:13
  wire            _T_1105;	// matmul/matmul-hw.mlir:16006:13
  wire            _T_1106;	// matmul/matmul-hw.mlir:16004:13
  wire            _T_1107;	// matmul/matmul-hw.mlir:16003:13
  wire [31:0]     _T_1108;	// matmul/matmul-hw.mlir:15994:13
  wire            _T_1109;	// matmul/matmul-hw.mlir:15993:13
  wire            _T_1110;	// matmul/matmul-hw.mlir:15976:13
  wire            _T_1111;	// matmul/matmul-hw.mlir:15974:13
  wire            _T_1112;	// matmul/matmul-hw.mlir:15973:13
  wire [31:0]     _T_1113;	// matmul/matmul-hw.mlir:15964:13
  wire            _T_1114;	// matmul/matmul-hw.mlir:15963:13
  wire            _T_1115;	// matmul/matmul-hw.mlir:15946:13
  wire            _T_1116;	// matmul/matmul-hw.mlir:15944:13
  wire            _T_1117;	// matmul/matmul-hw.mlir:15943:13
  wire [31:0]     _T_1118;	// matmul/matmul-hw.mlir:15934:13
  wire            _T_1119;	// matmul/matmul-hw.mlir:15933:13
  wire            _T_1120;	// matmul/matmul-hw.mlir:15916:13
  wire            _T_1121;	// matmul/matmul-hw.mlir:15914:13
  wire            _T_1122;	// matmul/matmul-hw.mlir:15913:13
  wire [31:0]     _T_1123;	// matmul/matmul-hw.mlir:15904:13
  wire            _T_1124;	// matmul/matmul-hw.mlir:15903:13
  wire            _T_1125;	// matmul/matmul-hw.mlir:15886:13
  wire            _T_1126;	// matmul/matmul-hw.mlir:15884:13
  wire            _T_1127;	// matmul/matmul-hw.mlir:15883:13
  wire [31:0]     _T_1128;	// matmul/matmul-hw.mlir:15882:13
  wire            _T_1129;	// matmul/matmul-hw.mlir:15881:13
  wire [31:0]     _T_1130;	// matmul/matmul-hw.mlir:15787:13
  wire            _T_1131;	// matmul/matmul-hw.mlir:15786:13
  wire [3:0]      _T_1132;	// matmul/matmul-hw.mlir:15785:13
  wire            _T_1133;	// matmul/matmul-hw.mlir:15784:13
  wire            _T_1134;	// matmul/matmul-hw.mlir:15768:13
  wire [31:0]     _T_1135;	// matmul/matmul-hw.mlir:15759:13
  wire            _T_1136;	// matmul/matmul-hw.mlir:15758:13
  wire            _T_1137;	// matmul/matmul-hw.mlir:15741:13
  wire            _T_1138;	// matmul/matmul-hw.mlir:15739:13
  wire            _T_1139;	// matmul/matmul-hw.mlir:15738:13
  wire [31:0]     _T_1140;	// matmul/matmul-hw.mlir:15729:13
  wire            _T_1141;	// matmul/matmul-hw.mlir:15728:13
  wire            _T_1142;	// matmul/matmul-hw.mlir:15711:13
  wire            _T_1143;	// matmul/matmul-hw.mlir:15709:13
  wire            _T_1144;	// matmul/matmul-hw.mlir:15708:13
  wire [31:0]     _T_1145;	// matmul/matmul-hw.mlir:15699:13
  wire            _T_1146;	// matmul/matmul-hw.mlir:15698:13
  wire            _T_1147;	// matmul/matmul-hw.mlir:15681:13
  wire            _T_1148;	// matmul/matmul-hw.mlir:15679:13
  wire            _T_1149;	// matmul/matmul-hw.mlir:15678:13
  wire [31:0]     _T_1150;	// matmul/matmul-hw.mlir:15669:13
  wire            _T_1151;	// matmul/matmul-hw.mlir:15668:13
  wire            _T_1152;	// matmul/matmul-hw.mlir:15651:13
  wire            _T_1153;	// matmul/matmul-hw.mlir:15649:13
  wire            _T_1154;	// matmul/matmul-hw.mlir:15648:13
  wire [31:0]     _T_1155;	// matmul/matmul-hw.mlir:15639:13
  wire            _T_1156;	// matmul/matmul-hw.mlir:15638:13
  wire            _T_1157;	// matmul/matmul-hw.mlir:15621:13
  wire            _T_1158;	// matmul/matmul-hw.mlir:15619:13
  wire            _T_1159;	// matmul/matmul-hw.mlir:15618:13
  wire [31:0]     _T_1160;	// matmul/matmul-hw.mlir:15609:13
  wire            _T_1161;	// matmul/matmul-hw.mlir:15608:13
  wire            _T_1162;	// matmul/matmul-hw.mlir:15591:13
  wire            _T_1163;	// matmul/matmul-hw.mlir:15589:13
  wire            _T_1164;	// matmul/matmul-hw.mlir:15588:13
  wire [31:0]     _T_1165;	// matmul/matmul-hw.mlir:15579:13
  wire            _T_1166;	// matmul/matmul-hw.mlir:15578:13
  wire            _T_1167;	// matmul/matmul-hw.mlir:15561:13
  wire            _T_1168;	// matmul/matmul-hw.mlir:15559:13
  wire            _T_1169;	// matmul/matmul-hw.mlir:15558:13
  wire [31:0]     _T_1170;	// matmul/matmul-hw.mlir:15549:13
  wire            _T_1171;	// matmul/matmul-hw.mlir:15548:13
  wire            _T_1172;	// matmul/matmul-hw.mlir:15531:13
  wire            _T_1173;	// matmul/matmul-hw.mlir:15529:13
  wire            _T_1174;	// matmul/matmul-hw.mlir:15528:13
  wire [31:0]     _T_1175;	// matmul/matmul-hw.mlir:15519:13
  wire            _T_1176;	// matmul/matmul-hw.mlir:15518:13
  wire            _T_1177;	// matmul/matmul-hw.mlir:15501:13
  wire            _T_1178;	// matmul/matmul-hw.mlir:15499:13
  wire            _T_1179;	// matmul/matmul-hw.mlir:15498:13
  wire [31:0]     _T_1180;	// matmul/matmul-hw.mlir:15489:13
  wire            _T_1181;	// matmul/matmul-hw.mlir:15488:13
  wire            _T_1182;	// matmul/matmul-hw.mlir:15471:13
  wire            _T_1183;	// matmul/matmul-hw.mlir:15469:13
  wire            _T_1184;	// matmul/matmul-hw.mlir:15468:13
  wire [31:0]     _T_1185;	// matmul/matmul-hw.mlir:15459:13
  wire            _T_1186;	// matmul/matmul-hw.mlir:15458:13
  wire            _T_1187;	// matmul/matmul-hw.mlir:15441:13
  wire            _T_1188;	// matmul/matmul-hw.mlir:15439:13
  wire            _T_1189;	// matmul/matmul-hw.mlir:15438:13
  wire [31:0]     _T_1190;	// matmul/matmul-hw.mlir:15429:13
  wire            _T_1191;	// matmul/matmul-hw.mlir:15428:13
  wire            _T_1192;	// matmul/matmul-hw.mlir:15411:13
  wire            _T_1193;	// matmul/matmul-hw.mlir:15409:13
  wire            _T_1194;	// matmul/matmul-hw.mlir:15408:13
  wire [31:0]     _T_1195;	// matmul/matmul-hw.mlir:15399:13
  wire            _T_1196;	// matmul/matmul-hw.mlir:15398:13
  wire            _T_1197;	// matmul/matmul-hw.mlir:15381:13
  wire            _T_1198;	// matmul/matmul-hw.mlir:15379:13
  wire            _T_1199;	// matmul/matmul-hw.mlir:15378:13
  wire [31:0]     _T_1200;	// matmul/matmul-hw.mlir:15369:13
  wire            _T_1201;	// matmul/matmul-hw.mlir:15368:13
  wire            _T_1202;	// matmul/matmul-hw.mlir:15351:13
  wire            _T_1203;	// matmul/matmul-hw.mlir:15349:13
  wire            _T_1204;	// matmul/matmul-hw.mlir:15348:13
  wire [31:0]     _T_1205;	// matmul/matmul-hw.mlir:15339:13
  wire            _T_1206;	// matmul/matmul-hw.mlir:15338:13
  wire            _T_1207;	// matmul/matmul-hw.mlir:15321:13
  wire            _T_1208;	// matmul/matmul-hw.mlir:15319:13
  wire            _T_1209;	// matmul/matmul-hw.mlir:15318:13
  wire [31:0]     _T_1210;	// matmul/matmul-hw.mlir:15309:13
  wire            _T_1211;	// matmul/matmul-hw.mlir:15308:13
  wire            _T_1212;	// matmul/matmul-hw.mlir:15291:13
  wire            _T_1213;	// matmul/matmul-hw.mlir:15289:13
  wire            _T_1214;	// matmul/matmul-hw.mlir:15288:13
  wire [31:0]     _T_1215;	// matmul/matmul-hw.mlir:15287:13
  wire            _T_1216;	// matmul/matmul-hw.mlir:15286:13
  wire [31:0]     _T_1217;	// matmul/matmul-hw.mlir:15192:13
  wire            _T_1218;	// matmul/matmul-hw.mlir:15191:13
  wire [3:0]      _T_1219;	// matmul/matmul-hw.mlir:15190:13
  wire            _T_1220;	// matmul/matmul-hw.mlir:15189:13
  wire            _T_1221;	// matmul/matmul-hw.mlir:15173:13
  wire [31:0]     _T_1222;	// matmul/matmul-hw.mlir:15164:13
  wire            _T_1223;	// matmul/matmul-hw.mlir:15163:13
  wire            _T_1224;	// matmul/matmul-hw.mlir:15146:13
  wire            _T_1225;	// matmul/matmul-hw.mlir:15144:13
  wire            _T_1226;	// matmul/matmul-hw.mlir:15143:13
  wire [31:0]     _T_1227;	// matmul/matmul-hw.mlir:15134:13
  wire            _T_1228;	// matmul/matmul-hw.mlir:15133:13
  wire            _T_1229;	// matmul/matmul-hw.mlir:15116:13
  wire            _T_1230;	// matmul/matmul-hw.mlir:15114:13
  wire            _T_1231;	// matmul/matmul-hw.mlir:15113:13
  wire [31:0]     _T_1232;	// matmul/matmul-hw.mlir:15104:13
  wire            _T_1233;	// matmul/matmul-hw.mlir:15103:13
  wire            _T_1234;	// matmul/matmul-hw.mlir:15086:13
  wire            _T_1235;	// matmul/matmul-hw.mlir:15084:13
  wire            _T_1236;	// matmul/matmul-hw.mlir:15083:13
  wire [31:0]     _T_1237;	// matmul/matmul-hw.mlir:15074:13
  wire            _T_1238;	// matmul/matmul-hw.mlir:15073:13
  wire            _T_1239;	// matmul/matmul-hw.mlir:15056:13
  wire            _T_1240;	// matmul/matmul-hw.mlir:15054:13
  wire            _T_1241;	// matmul/matmul-hw.mlir:15053:13
  wire [31:0]     _T_1242;	// matmul/matmul-hw.mlir:15044:13
  wire            _T_1243;	// matmul/matmul-hw.mlir:15043:13
  wire            _T_1244;	// matmul/matmul-hw.mlir:15026:13
  wire            _T_1245;	// matmul/matmul-hw.mlir:15024:13
  wire            _T_1246;	// matmul/matmul-hw.mlir:15023:13
  wire [31:0]     _T_1247;	// matmul/matmul-hw.mlir:15014:13
  wire            _T_1248;	// matmul/matmul-hw.mlir:15013:13
  wire            _T_1249;	// matmul/matmul-hw.mlir:14996:13
  wire            _T_1250;	// matmul/matmul-hw.mlir:14994:13
  wire            _T_1251;	// matmul/matmul-hw.mlir:14993:13
  wire [31:0]     _T_1252;	// matmul/matmul-hw.mlir:14984:13
  wire            _T_1253;	// matmul/matmul-hw.mlir:14983:13
  wire            _T_1254;	// matmul/matmul-hw.mlir:14966:13
  wire            _T_1255;	// matmul/matmul-hw.mlir:14964:13
  wire            _T_1256;	// matmul/matmul-hw.mlir:14963:13
  wire [31:0]     _T_1257;	// matmul/matmul-hw.mlir:14954:13
  wire            _T_1258;	// matmul/matmul-hw.mlir:14953:13
  wire            _T_1259;	// matmul/matmul-hw.mlir:14936:13
  wire            _T_1260;	// matmul/matmul-hw.mlir:14934:13
  wire            _T_1261;	// matmul/matmul-hw.mlir:14933:13
  wire [31:0]     _T_1262;	// matmul/matmul-hw.mlir:14924:13
  wire            _T_1263;	// matmul/matmul-hw.mlir:14923:13
  wire            _T_1264;	// matmul/matmul-hw.mlir:14906:13
  wire            _T_1265;	// matmul/matmul-hw.mlir:14904:13
  wire            _T_1266;	// matmul/matmul-hw.mlir:14903:13
  wire [31:0]     _T_1267;	// matmul/matmul-hw.mlir:14894:13
  wire            _T_1268;	// matmul/matmul-hw.mlir:14893:13
  wire            _T_1269;	// matmul/matmul-hw.mlir:14876:13
  wire            _T_1270;	// matmul/matmul-hw.mlir:14874:13
  wire            _T_1271;	// matmul/matmul-hw.mlir:14873:13
  wire [31:0]     _T_1272;	// matmul/matmul-hw.mlir:14864:13
  wire            _T_1273;	// matmul/matmul-hw.mlir:14863:13
  wire            _T_1274;	// matmul/matmul-hw.mlir:14846:13
  wire            _T_1275;	// matmul/matmul-hw.mlir:14844:13
  wire            _T_1276;	// matmul/matmul-hw.mlir:14843:13
  wire [31:0]     _T_1277;	// matmul/matmul-hw.mlir:14834:13
  wire            _T_1278;	// matmul/matmul-hw.mlir:14833:13
  wire            _T_1279;	// matmul/matmul-hw.mlir:14816:13
  wire            _T_1280;	// matmul/matmul-hw.mlir:14814:13
  wire            _T_1281;	// matmul/matmul-hw.mlir:14813:13
  wire [31:0]     _T_1282;	// matmul/matmul-hw.mlir:14804:13
  wire            _T_1283;	// matmul/matmul-hw.mlir:14803:13
  wire            _T_1284;	// matmul/matmul-hw.mlir:14786:13
  wire            _T_1285;	// matmul/matmul-hw.mlir:14784:13
  wire            _T_1286;	// matmul/matmul-hw.mlir:14783:13
  wire [31:0]     _T_1287;	// matmul/matmul-hw.mlir:14774:13
  wire            _T_1288;	// matmul/matmul-hw.mlir:14773:13
  wire            _T_1289;	// matmul/matmul-hw.mlir:14756:13
  wire            _T_1290;	// matmul/matmul-hw.mlir:14754:13
  wire            _T_1291;	// matmul/matmul-hw.mlir:14753:13
  wire [31:0]     _T_1292;	// matmul/matmul-hw.mlir:14744:13
  wire            _T_1293;	// matmul/matmul-hw.mlir:14743:13
  wire            _T_1294;	// matmul/matmul-hw.mlir:14726:13
  wire            _T_1295;	// matmul/matmul-hw.mlir:14724:13
  wire            _T_1296;	// matmul/matmul-hw.mlir:14723:13
  wire [31:0]     _T_1297;	// matmul/matmul-hw.mlir:14714:13
  wire            _T_1298;	// matmul/matmul-hw.mlir:14713:13
  wire            _T_1299;	// matmul/matmul-hw.mlir:14696:13
  wire            _T_1300;	// matmul/matmul-hw.mlir:14694:13
  wire            _T_1301;	// matmul/matmul-hw.mlir:14693:13
  wire [31:0]     _T_1302;	// matmul/matmul-hw.mlir:14692:13
  wire            _T_1303;	// matmul/matmul-hw.mlir:14691:13
  wire [31:0]     _T_1304;	// matmul/matmul-hw.mlir:14597:13
  wire            _T_1305;	// matmul/matmul-hw.mlir:14596:13
  wire [3:0]      _T_1306;	// matmul/matmul-hw.mlir:14595:13
  wire            _T_1307;	// matmul/matmul-hw.mlir:14594:13
  wire            _T_1308;	// matmul/matmul-hw.mlir:14578:13
  wire [31:0]     _T_1309;	// matmul/matmul-hw.mlir:14577:13
  wire            _T_1310;	// matmul/matmul-hw.mlir:14576:13
  wire            _T_1311;	// matmul/matmul-hw.mlir:14559:13
  wire            _T_1312;	// matmul/matmul-hw.mlir:14557:13
  wire            _T_1313;	// matmul/matmul-hw.mlir:14556:13
  wire [31:0]     _T_1314;	// matmul/matmul-hw.mlir:14555:13
  wire            _T_1315;	// matmul/matmul-hw.mlir:14554:13
  wire            _T_1316;	// matmul/matmul-hw.mlir:14537:13
  wire            _T_1317;	// matmul/matmul-hw.mlir:14535:13
  wire            _T_1318;	// matmul/matmul-hw.mlir:14534:13
  wire [31:0]     _T_1319;	// matmul/matmul-hw.mlir:14533:13
  wire            _T_1320;	// matmul/matmul-hw.mlir:14532:13
  wire            _T_1321;	// matmul/matmul-hw.mlir:14515:13
  wire            _T_1322;	// matmul/matmul-hw.mlir:14513:13
  wire            _T_1323;	// matmul/matmul-hw.mlir:14512:13
  wire [31:0]     _T_1324;	// matmul/matmul-hw.mlir:14511:13
  wire            _T_1325;	// matmul/matmul-hw.mlir:14510:13
  wire            _T_1326;	// matmul/matmul-hw.mlir:14493:13
  wire            _T_1327;	// matmul/matmul-hw.mlir:14491:13
  wire            _T_1328;	// matmul/matmul-hw.mlir:14490:13
  wire [31:0]     _T_1329;	// matmul/matmul-hw.mlir:14489:13
  wire            _T_1330;	// matmul/matmul-hw.mlir:14488:13
  wire            _T_1331;	// matmul/matmul-hw.mlir:14471:13
  wire            _T_1332;	// matmul/matmul-hw.mlir:14469:13
  wire            _T_1333;	// matmul/matmul-hw.mlir:14468:13
  wire [31:0]     _T_1334;	// matmul/matmul-hw.mlir:14467:13
  wire            _T_1335;	// matmul/matmul-hw.mlir:14466:13
  wire            _T_1336;	// matmul/matmul-hw.mlir:14449:13
  wire            _T_1337;	// matmul/matmul-hw.mlir:14447:13
  wire            _T_1338;	// matmul/matmul-hw.mlir:14446:13
  wire [31:0]     _T_1339;	// matmul/matmul-hw.mlir:14445:13
  wire            _T_1340;	// matmul/matmul-hw.mlir:14444:13
  wire            _T_1341;	// matmul/matmul-hw.mlir:14427:13
  wire            _T_1342;	// matmul/matmul-hw.mlir:14425:13
  wire            _T_1343;	// matmul/matmul-hw.mlir:14424:13
  wire [31:0]     _T_1344;	// matmul/matmul-hw.mlir:14423:13
  wire            _T_1345;	// matmul/matmul-hw.mlir:14422:13
  wire            _T_1346;	// matmul/matmul-hw.mlir:14405:13
  wire            _T_1347;	// matmul/matmul-hw.mlir:14403:13
  wire            _T_1348;	// matmul/matmul-hw.mlir:14402:13
  wire [31:0]     _T_1349;	// matmul/matmul-hw.mlir:14401:13
  wire            _T_1350;	// matmul/matmul-hw.mlir:14400:13
  wire            _T_1351;	// matmul/matmul-hw.mlir:14383:13
  wire            _T_1352;	// matmul/matmul-hw.mlir:14381:13
  wire            _T_1353;	// matmul/matmul-hw.mlir:14380:13
  wire [31:0]     _T_1354;	// matmul/matmul-hw.mlir:14379:13
  wire            _T_1355;	// matmul/matmul-hw.mlir:14378:13
  wire            _T_1356;	// matmul/matmul-hw.mlir:14361:13
  wire            _T_1357;	// matmul/matmul-hw.mlir:14359:13
  wire            _T_1358;	// matmul/matmul-hw.mlir:14358:13
  wire [31:0]     _T_1359;	// matmul/matmul-hw.mlir:14357:13
  wire            _T_1360;	// matmul/matmul-hw.mlir:14356:13
  wire            _T_1361;	// matmul/matmul-hw.mlir:14339:13
  wire            _T_1362;	// matmul/matmul-hw.mlir:14337:13
  wire            _T_1363;	// matmul/matmul-hw.mlir:14336:13
  wire [31:0]     _T_1364;	// matmul/matmul-hw.mlir:14335:13
  wire            _T_1365;	// matmul/matmul-hw.mlir:14334:13
  wire            _T_1366;	// matmul/matmul-hw.mlir:14317:13
  wire            _T_1367;	// matmul/matmul-hw.mlir:14315:13
  wire            _T_1368;	// matmul/matmul-hw.mlir:14314:13
  wire [31:0]     _T_1369;	// matmul/matmul-hw.mlir:14313:13
  wire            _T_1370;	// matmul/matmul-hw.mlir:14312:13
  wire            _T_1371;	// matmul/matmul-hw.mlir:14295:13
  wire            _T_1372;	// matmul/matmul-hw.mlir:14293:13
  wire            _T_1373;	// matmul/matmul-hw.mlir:14292:13
  wire [31:0]     _T_1374;	// matmul/matmul-hw.mlir:14291:13
  wire            _T_1375;	// matmul/matmul-hw.mlir:14290:13
  wire            _T_1376;	// matmul/matmul-hw.mlir:14273:13
  wire            _T_1377;	// matmul/matmul-hw.mlir:14271:13
  wire            _T_1378;	// matmul/matmul-hw.mlir:14270:13
  wire [31:0]     _T_1379;	// matmul/matmul-hw.mlir:14269:13
  wire            _T_1380;	// matmul/matmul-hw.mlir:14268:13
  wire            _T_1381;	// matmul/matmul-hw.mlir:14251:13
  wire            _T_1382;	// matmul/matmul-hw.mlir:14249:13
  wire            _T_1383;	// matmul/matmul-hw.mlir:14248:13
  wire [31:0]     _T_1384;	// matmul/matmul-hw.mlir:14247:13
  wire            _T_1385;	// matmul/matmul-hw.mlir:14246:13
  wire            _T_1386;	// matmul/matmul-hw.mlir:14229:13
  wire            _T_1387;	// matmul/matmul-hw.mlir:14227:13
  wire            _T_1388;	// matmul/matmul-hw.mlir:14226:13
  wire [31:0]     _T_1389;	// matmul/matmul-hw.mlir:14225:13
  wire            _T_1390;	// matmul/matmul-hw.mlir:14224:13
  wire [31:0]     _T_1391;	// matmul/matmul-hw.mlir:14138:13
  wire            _T_1392;	// matmul/matmul-hw.mlir:14137:13
  wire            _T_1393;	// matmul/matmul-hw.mlir:14136:13
  wire [31:0]     _T_1394;	// matmul/matmul-hw.mlir:14120:13
  wire            _T_1395;	// matmul/matmul-hw.mlir:14119:13
  wire            _T_1396;	// matmul/matmul-hw.mlir:14118:13
  wire [31:0]     _T_1397;	// matmul/matmul-hw.mlir:14117:13
  wire            _T_1398;	// matmul/matmul-hw.mlir:14116:13
  wire            _T_1399;	// matmul/matmul-hw.mlir:14115:13
  wire [31:0]     _T_1400;	// matmul/matmul-hw.mlir:14114:13
  wire            _T_1401;	// matmul/matmul-hw.mlir:14113:13
  wire            _T_1402;	// matmul/matmul-hw.mlir:14112:13
  wire [31:0]     _T_1403;	// matmul/matmul-hw.mlir:14111:13
  wire            _T_1404;	// matmul/matmul-hw.mlir:14110:13
  wire            _T_1405;	// matmul/matmul-hw.mlir:14109:13
  wire [31:0]     _T_1406;	// matmul/matmul-hw.mlir:14108:13
  wire            _T_1407;	// matmul/matmul-hw.mlir:14107:13
  wire            _T_1408;	// matmul/matmul-hw.mlir:14106:13
  wire [31:0]     _T_1409;	// matmul/matmul-hw.mlir:14105:13
  wire            _T_1410;	// matmul/matmul-hw.mlir:14104:13
  wire            _T_1411;	// matmul/matmul-hw.mlir:14103:13
  wire [31:0]     _T_1412;	// matmul/matmul-hw.mlir:14102:13
  wire            _T_1413;	// matmul/matmul-hw.mlir:14101:13
  wire            _T_1414;	// matmul/matmul-hw.mlir:14100:13
  wire [31:0]     _T_1415;	// matmul/matmul-hw.mlir:14099:13
  wire            _T_1416;	// matmul/matmul-hw.mlir:14098:13
  wire            _T_1417;	// matmul/matmul-hw.mlir:14097:13
  wire [31:0]     _T_1418;	// matmul/matmul-hw.mlir:14096:13
  wire            _T_1419;	// matmul/matmul-hw.mlir:14095:13
  wire            _T_1420;	// matmul/matmul-hw.mlir:14094:13
  wire [31:0]     _T_1421;	// matmul/matmul-hw.mlir:14093:13
  wire            _T_1422;	// matmul/matmul-hw.mlir:14092:13
  wire            _T_1423;	// matmul/matmul-hw.mlir:14091:13
  wire [31:0]     _T_1424;	// matmul/matmul-hw.mlir:14090:13
  wire            _T_1425;	// matmul/matmul-hw.mlir:14089:13
  wire            _T_1426;	// matmul/matmul-hw.mlir:14088:13
  wire [31:0]     _T_1427;	// matmul/matmul-hw.mlir:14087:13
  wire            _T_1428;	// matmul/matmul-hw.mlir:14086:13
  wire            _T_1429;	// matmul/matmul-hw.mlir:14085:13
  wire [31:0]     _T_1430;	// matmul/matmul-hw.mlir:14084:13
  wire            _T_1431;	// matmul/matmul-hw.mlir:14083:13
  wire            _T_1432;	// matmul/matmul-hw.mlir:14082:13
  wire [31:0]     _T_1433;	// matmul/matmul-hw.mlir:14081:13
  wire            _T_1434;	// matmul/matmul-hw.mlir:14080:13
  wire            _T_1435;	// matmul/matmul-hw.mlir:14079:13
  wire [31:0]     _T_1436;	// matmul/matmul-hw.mlir:14078:13
  wire            _T_1437;	// matmul/matmul-hw.mlir:14077:13
  wire            _T_1438;	// matmul/matmul-hw.mlir:14076:13
  wire [31:0]     _T_1439;	// matmul/matmul-hw.mlir:14075:13
  wire            _T_1440;	// matmul/matmul-hw.mlir:14074:13
  wire            _T_1441;	// matmul/matmul-hw.mlir:14073:13
  wire [31:0]     _T_1442;	// matmul/matmul-hw.mlir:14057:13
  wire            _T_1443;	// matmul/matmul-hw.mlir:14056:13
  wire            _T_1444;	// matmul/matmul-hw.mlir:14055:13
  wire [31:0]     _T_1445;	// matmul/matmul-hw.mlir:14054:13
  wire            _T_1446;	// matmul/matmul-hw.mlir:14053:13
  wire            _T_1447;	// matmul/matmul-hw.mlir:14052:13
  wire [31:0]     _T_1448;	// matmul/matmul-hw.mlir:14051:13
  wire            _T_1449;	// matmul/matmul-hw.mlir:14050:13
  wire            _T_1450;	// matmul/matmul-hw.mlir:14049:13
  wire [31:0]     _T_1451;	// matmul/matmul-hw.mlir:14048:13
  wire            _T_1452;	// matmul/matmul-hw.mlir:14047:13
  wire            _T_1453;	// matmul/matmul-hw.mlir:14046:13
  wire [31:0]     _T_1454;	// matmul/matmul-hw.mlir:14045:13
  wire            _T_1455;	// matmul/matmul-hw.mlir:14044:13
  wire            _T_1456;	// matmul/matmul-hw.mlir:14043:13
  wire [31:0]     _T_1457;	// matmul/matmul-hw.mlir:14042:13
  wire            _T_1458;	// matmul/matmul-hw.mlir:14041:13
  wire            _T_1459;	// matmul/matmul-hw.mlir:14040:13
  wire [31:0]     _T_1460;	// matmul/matmul-hw.mlir:14039:13
  wire            _T_1461;	// matmul/matmul-hw.mlir:14038:13
  wire            _T_1462;	// matmul/matmul-hw.mlir:14037:13
  wire [31:0]     _T_1463;	// matmul/matmul-hw.mlir:14036:13
  wire            _T_1464;	// matmul/matmul-hw.mlir:14035:13
  wire            _T_1465;	// matmul/matmul-hw.mlir:14034:13
  wire [31:0]     _T_1466;	// matmul/matmul-hw.mlir:14033:13
  wire            _T_1467;	// matmul/matmul-hw.mlir:14032:13
  wire            _T_1468;	// matmul/matmul-hw.mlir:14031:13
  wire [31:0]     _T_1469;	// matmul/matmul-hw.mlir:14030:13
  wire            _T_1470;	// matmul/matmul-hw.mlir:14029:13
  wire            _T_1471;	// matmul/matmul-hw.mlir:14028:13
  wire [31:0]     _T_1472;	// matmul/matmul-hw.mlir:14027:13
  wire            _T_1473;	// matmul/matmul-hw.mlir:14026:13
  wire            _T_1474;	// matmul/matmul-hw.mlir:14025:13
  wire [31:0]     _T_1475;	// matmul/matmul-hw.mlir:14024:13
  wire            _T_1476;	// matmul/matmul-hw.mlir:14023:13
  wire            _T_1477;	// matmul/matmul-hw.mlir:14022:13
  wire [31:0]     _T_1478;	// matmul/matmul-hw.mlir:14021:13
  wire            _T_1479;	// matmul/matmul-hw.mlir:14020:13
  wire            _T_1480;	// matmul/matmul-hw.mlir:14019:13
  wire [31:0]     _T_1481;	// matmul/matmul-hw.mlir:14018:13
  wire            _T_1482;	// matmul/matmul-hw.mlir:14017:13
  wire            _T_1483;	// matmul/matmul-hw.mlir:14016:13
  wire [31:0]     _T_1484;	// matmul/matmul-hw.mlir:14015:13
  wire            _T_1485;	// matmul/matmul-hw.mlir:14014:13
  wire            _T_1486;	// matmul/matmul-hw.mlir:14013:13
  wire [31:0]     _T_1487;	// matmul/matmul-hw.mlir:14012:13
  wire            _T_1488;	// matmul/matmul-hw.mlir:14011:13
  wire            _T_1489;	// matmul/matmul-hw.mlir:14010:13
  wire [31:0]     _T_1490;	// matmul/matmul-hw.mlir:13994:13
  wire            _T_1491;	// matmul/matmul-hw.mlir:13993:13
  wire            _T_1492;	// matmul/matmul-hw.mlir:13992:13
  wire [31:0]     _T_1493;	// matmul/matmul-hw.mlir:13991:13
  wire            _T_1494;	// matmul/matmul-hw.mlir:13990:13
  wire            _T_1495;	// matmul/matmul-hw.mlir:13989:13
  wire [31:0]     _T_1496;	// matmul/matmul-hw.mlir:13988:13
  wire            _T_1497;	// matmul/matmul-hw.mlir:13987:13
  wire            _T_1498;	// matmul/matmul-hw.mlir:13986:13
  wire [31:0]     _T_1499;	// matmul/matmul-hw.mlir:13985:13
  wire            _T_1500;	// matmul/matmul-hw.mlir:13984:13
  wire            _T_1501;	// matmul/matmul-hw.mlir:13983:13
  wire [31:0]     _T_1502;	// matmul/matmul-hw.mlir:13982:13
  wire            _T_1503;	// matmul/matmul-hw.mlir:13981:13
  wire            _T_1504;	// matmul/matmul-hw.mlir:13980:13
  wire [31:0]     _T_1505;	// matmul/matmul-hw.mlir:13979:13
  wire            _T_1506;	// matmul/matmul-hw.mlir:13978:13
  wire            _T_1507;	// matmul/matmul-hw.mlir:13977:13
  wire [31:0]     _T_1508;	// matmul/matmul-hw.mlir:13976:13
  wire            _T_1509;	// matmul/matmul-hw.mlir:13975:13
  wire            _T_1510;	// matmul/matmul-hw.mlir:13974:13
  wire [31:0]     _T_1511;	// matmul/matmul-hw.mlir:13973:13
  wire            _T_1512;	// matmul/matmul-hw.mlir:13972:13
  wire            _T_1513;	// matmul/matmul-hw.mlir:13971:13
  wire [31:0]     _T_1514;	// matmul/matmul-hw.mlir:13970:13
  wire            _T_1515;	// matmul/matmul-hw.mlir:13969:13
  wire            _T_1516;	// matmul/matmul-hw.mlir:13968:13
  wire [31:0]     _T_1517;	// matmul/matmul-hw.mlir:13967:13
  wire            _T_1518;	// matmul/matmul-hw.mlir:13966:13
  wire            _T_1519;	// matmul/matmul-hw.mlir:13965:13
  wire [31:0]     _T_1520;	// matmul/matmul-hw.mlir:13964:13
  wire            _T_1521;	// matmul/matmul-hw.mlir:13963:13
  wire            _T_1522;	// matmul/matmul-hw.mlir:13962:13
  wire [31:0]     _T_1523;	// matmul/matmul-hw.mlir:13961:13
  wire            _T_1524;	// matmul/matmul-hw.mlir:13960:13
  wire            _T_1525;	// matmul/matmul-hw.mlir:13959:13
  wire [31:0]     _T_1526;	// matmul/matmul-hw.mlir:13958:13
  wire            _T_1527;	// matmul/matmul-hw.mlir:13957:13
  wire            _T_1528;	// matmul/matmul-hw.mlir:13956:13
  wire [31:0]     _T_1529;	// matmul/matmul-hw.mlir:13955:13
  wire            _T_1530;	// matmul/matmul-hw.mlir:13954:13
  wire            _T_1531;	// matmul/matmul-hw.mlir:13953:13
  wire [31:0]     _T_1532;	// matmul/matmul-hw.mlir:13952:13
  wire            _T_1533;	// matmul/matmul-hw.mlir:13951:13
  wire            _T_1534;	// matmul/matmul-hw.mlir:13950:13
  wire [31:0]     _T_1535;	// matmul/matmul-hw.mlir:13949:13
  wire            _T_1536;	// matmul/matmul-hw.mlir:13948:13
  wire            _T_1537;	// matmul/matmul-hw.mlir:13947:13
  wire [31:0]     _T_1538;	// matmul/matmul-hw.mlir:13931:13
  wire            _T_1539;	// matmul/matmul-hw.mlir:13930:13
  wire            _T_1540;	// matmul/matmul-hw.mlir:13929:13
  wire [31:0]     _T_1541;	// matmul/matmul-hw.mlir:13928:13
  wire            _T_1542;	// matmul/matmul-hw.mlir:13927:13
  wire            _T_1543;	// matmul/matmul-hw.mlir:13926:13
  wire [31:0]     _T_1544;	// matmul/matmul-hw.mlir:13925:13
  wire            _T_1545;	// matmul/matmul-hw.mlir:13924:13
  wire            _T_1546;	// matmul/matmul-hw.mlir:13923:13
  wire [31:0]     _T_1547;	// matmul/matmul-hw.mlir:13922:13
  wire            _T_1548;	// matmul/matmul-hw.mlir:13921:13
  wire            _T_1549;	// matmul/matmul-hw.mlir:13920:13
  wire [31:0]     _T_1550;	// matmul/matmul-hw.mlir:13919:13
  wire            _T_1551;	// matmul/matmul-hw.mlir:13918:13
  wire            _T_1552;	// matmul/matmul-hw.mlir:13917:13
  wire [31:0]     _T_1553;	// matmul/matmul-hw.mlir:13916:13
  wire            _T_1554;	// matmul/matmul-hw.mlir:13915:13
  wire            _T_1555;	// matmul/matmul-hw.mlir:13914:13
  wire [31:0]     _T_1556;	// matmul/matmul-hw.mlir:13913:13
  wire            _T_1557;	// matmul/matmul-hw.mlir:13912:13
  wire            _T_1558;	// matmul/matmul-hw.mlir:13911:13
  wire [31:0]     _T_1559;	// matmul/matmul-hw.mlir:13910:13
  wire            _T_1560;	// matmul/matmul-hw.mlir:13909:13
  wire            _T_1561;	// matmul/matmul-hw.mlir:13908:13
  wire [31:0]     _T_1562;	// matmul/matmul-hw.mlir:13907:13
  wire            _T_1563;	// matmul/matmul-hw.mlir:13906:13
  wire            _T_1564;	// matmul/matmul-hw.mlir:13905:13
  wire [31:0]     _T_1565;	// matmul/matmul-hw.mlir:13904:13
  wire            _T_1566;	// matmul/matmul-hw.mlir:13903:13
  wire            _T_1567;	// matmul/matmul-hw.mlir:13902:13
  wire [31:0]     _T_1568;	// matmul/matmul-hw.mlir:13901:13
  wire            _T_1569;	// matmul/matmul-hw.mlir:13900:13
  wire            _T_1570;	// matmul/matmul-hw.mlir:13899:13
  wire [31:0]     _T_1571;	// matmul/matmul-hw.mlir:13898:13
  wire            _T_1572;	// matmul/matmul-hw.mlir:13897:13
  wire            _T_1573;	// matmul/matmul-hw.mlir:13896:13
  wire [31:0]     _T_1574;	// matmul/matmul-hw.mlir:13895:13
  wire            _T_1575;	// matmul/matmul-hw.mlir:13894:13
  wire            _T_1576;	// matmul/matmul-hw.mlir:13893:13
  wire [31:0]     _T_1577;	// matmul/matmul-hw.mlir:13892:13
  wire            _T_1578;	// matmul/matmul-hw.mlir:13891:13
  wire            _T_1579;	// matmul/matmul-hw.mlir:13890:13
  wire [31:0]     _T_1580;	// matmul/matmul-hw.mlir:13889:13
  wire            _T_1581;	// matmul/matmul-hw.mlir:13888:13
  wire            _T_1582;	// matmul/matmul-hw.mlir:13887:13
  wire [31:0]     _T_1583;	// matmul/matmul-hw.mlir:13886:13
  wire            _T_1584;	// matmul/matmul-hw.mlir:13885:13
  wire            _T_1585;	// matmul/matmul-hw.mlir:13884:13
  wire [31:0]     _T_1586;	// matmul/matmul-hw.mlir:13868:13
  wire            _T_1587;	// matmul/matmul-hw.mlir:13867:13
  wire            _T_1588;	// matmul/matmul-hw.mlir:13866:13
  wire [31:0]     _T_1589;	// matmul/matmul-hw.mlir:13865:13
  wire            _T_1590;	// matmul/matmul-hw.mlir:13864:13
  wire            _T_1591;	// matmul/matmul-hw.mlir:13863:13
  wire [31:0]     _T_1592;	// matmul/matmul-hw.mlir:13862:13
  wire            _T_1593;	// matmul/matmul-hw.mlir:13861:13
  wire            _T_1594;	// matmul/matmul-hw.mlir:13860:13
  wire [31:0]     _T_1595;	// matmul/matmul-hw.mlir:13859:13
  wire            _T_1596;	// matmul/matmul-hw.mlir:13858:13
  wire            _T_1597;	// matmul/matmul-hw.mlir:13857:13
  wire [31:0]     _T_1598;	// matmul/matmul-hw.mlir:13856:13
  wire            _T_1599;	// matmul/matmul-hw.mlir:13855:13
  wire            _T_1600;	// matmul/matmul-hw.mlir:13854:13
  wire [31:0]     _T_1601;	// matmul/matmul-hw.mlir:13853:13
  wire            _T_1602;	// matmul/matmul-hw.mlir:13852:13
  wire            _T_1603;	// matmul/matmul-hw.mlir:13851:13
  wire [31:0]     _T_1604;	// matmul/matmul-hw.mlir:13850:13
  wire            _T_1605;	// matmul/matmul-hw.mlir:13849:13
  wire            _T_1606;	// matmul/matmul-hw.mlir:13848:13
  wire [31:0]     _T_1607;	// matmul/matmul-hw.mlir:13847:13
  wire            _T_1608;	// matmul/matmul-hw.mlir:13846:13
  wire            _T_1609;	// matmul/matmul-hw.mlir:13845:13
  wire [31:0]     _T_1610;	// matmul/matmul-hw.mlir:13844:13
  wire            _T_1611;	// matmul/matmul-hw.mlir:13843:13
  wire            _T_1612;	// matmul/matmul-hw.mlir:13842:13
  wire [31:0]     _T_1613;	// matmul/matmul-hw.mlir:13841:13
  wire            _T_1614;	// matmul/matmul-hw.mlir:13840:13
  wire            _T_1615;	// matmul/matmul-hw.mlir:13839:13
  wire [31:0]     _T_1616;	// matmul/matmul-hw.mlir:13838:13
  wire            _T_1617;	// matmul/matmul-hw.mlir:13837:13
  wire            _T_1618;	// matmul/matmul-hw.mlir:13836:13
  wire [31:0]     _T_1619;	// matmul/matmul-hw.mlir:13835:13
  wire            _T_1620;	// matmul/matmul-hw.mlir:13834:13
  wire            _T_1621;	// matmul/matmul-hw.mlir:13833:13
  wire [31:0]     _T_1622;	// matmul/matmul-hw.mlir:13832:13
  wire            _T_1623;	// matmul/matmul-hw.mlir:13831:13
  wire            _T_1624;	// matmul/matmul-hw.mlir:13830:13
  wire [31:0]     _T_1625;	// matmul/matmul-hw.mlir:13829:13
  wire            _T_1626;	// matmul/matmul-hw.mlir:13828:13
  wire            _T_1627;	// matmul/matmul-hw.mlir:13827:13
  wire [31:0]     _T_1628;	// matmul/matmul-hw.mlir:13826:13
  wire            _T_1629;	// matmul/matmul-hw.mlir:13825:13
  wire            _T_1630;	// matmul/matmul-hw.mlir:13824:13
  wire [31:0]     _T_1631;	// matmul/matmul-hw.mlir:13823:13
  wire            _T_1632;	// matmul/matmul-hw.mlir:13822:13
  wire            _T_1633;	// matmul/matmul-hw.mlir:13821:13
  wire [31:0]     _T_1634;	// matmul/matmul-hw.mlir:13805:13
  wire            _T_1635;	// matmul/matmul-hw.mlir:13804:13
  wire            _T_1636;	// matmul/matmul-hw.mlir:13803:13
  wire [31:0]     _T_1637;	// matmul/matmul-hw.mlir:13802:13
  wire            _T_1638;	// matmul/matmul-hw.mlir:13801:13
  wire            _T_1639;	// matmul/matmul-hw.mlir:13800:13
  wire [31:0]     _T_1640;	// matmul/matmul-hw.mlir:13799:13
  wire            _T_1641;	// matmul/matmul-hw.mlir:13798:13
  wire            _T_1642;	// matmul/matmul-hw.mlir:13797:13
  wire [31:0]     _T_1643;	// matmul/matmul-hw.mlir:13796:13
  wire            _T_1644;	// matmul/matmul-hw.mlir:13795:13
  wire            _T_1645;	// matmul/matmul-hw.mlir:13794:13
  wire [31:0]     _T_1646;	// matmul/matmul-hw.mlir:13793:13
  wire            _T_1647;	// matmul/matmul-hw.mlir:13792:13
  wire            _T_1648;	// matmul/matmul-hw.mlir:13791:13
  wire [31:0]     _T_1649;	// matmul/matmul-hw.mlir:13790:13
  wire            _T_1650;	// matmul/matmul-hw.mlir:13789:13
  wire            _T_1651;	// matmul/matmul-hw.mlir:13788:13
  wire [31:0]     _T_1652;	// matmul/matmul-hw.mlir:13787:13
  wire            _T_1653;	// matmul/matmul-hw.mlir:13786:13
  wire            _T_1654;	// matmul/matmul-hw.mlir:13785:13
  wire [31:0]     _T_1655;	// matmul/matmul-hw.mlir:13784:13
  wire            _T_1656;	// matmul/matmul-hw.mlir:13783:13
  wire            _T_1657;	// matmul/matmul-hw.mlir:13782:13
  wire [31:0]     _T_1658;	// matmul/matmul-hw.mlir:13781:13
  wire            _T_1659;	// matmul/matmul-hw.mlir:13780:13
  wire            _T_1660;	// matmul/matmul-hw.mlir:13779:13
  wire [31:0]     _T_1661;	// matmul/matmul-hw.mlir:13778:13
  wire            _T_1662;	// matmul/matmul-hw.mlir:13777:13
  wire            _T_1663;	// matmul/matmul-hw.mlir:13776:13
  wire [31:0]     _T_1664;	// matmul/matmul-hw.mlir:13775:13
  wire            _T_1665;	// matmul/matmul-hw.mlir:13774:13
  wire            _T_1666;	// matmul/matmul-hw.mlir:13773:13
  wire [31:0]     _T_1667;	// matmul/matmul-hw.mlir:13772:13
  wire            _T_1668;	// matmul/matmul-hw.mlir:13771:13
  wire            _T_1669;	// matmul/matmul-hw.mlir:13770:13
  wire [31:0]     _T_1670;	// matmul/matmul-hw.mlir:13769:13
  wire            _T_1671;	// matmul/matmul-hw.mlir:13768:13
  wire            _T_1672;	// matmul/matmul-hw.mlir:13767:13
  wire [31:0]     _T_1673;	// matmul/matmul-hw.mlir:13766:13
  wire            _T_1674;	// matmul/matmul-hw.mlir:13765:13
  wire            _T_1675;	// matmul/matmul-hw.mlir:13764:13
  wire [31:0]     _T_1676;	// matmul/matmul-hw.mlir:13763:13
  wire            _T_1677;	// matmul/matmul-hw.mlir:13762:13
  wire            _T_1678;	// matmul/matmul-hw.mlir:13761:13
  wire [31:0]     _T_1679;	// matmul/matmul-hw.mlir:13760:13
  wire            _T_1680;	// matmul/matmul-hw.mlir:13759:13
  wire            _T_1681;	// matmul/matmul-hw.mlir:13758:13
  wire [31:0]     _T_1682;	// matmul/matmul-hw.mlir:13742:13
  wire            _T_1683;	// matmul/matmul-hw.mlir:13741:13
  wire            _T_1684;	// matmul/matmul-hw.mlir:13740:13
  wire [31:0]     _T_1685;	// matmul/matmul-hw.mlir:13739:13
  wire            _T_1686;	// matmul/matmul-hw.mlir:13738:13
  wire            _T_1687;	// matmul/matmul-hw.mlir:13737:13
  wire [31:0]     _T_1688;	// matmul/matmul-hw.mlir:13736:13
  wire            _T_1689;	// matmul/matmul-hw.mlir:13735:13
  wire            _T_1690;	// matmul/matmul-hw.mlir:13734:13
  wire [31:0]     _T_1691;	// matmul/matmul-hw.mlir:13733:13
  wire            _T_1692;	// matmul/matmul-hw.mlir:13732:13
  wire            _T_1693;	// matmul/matmul-hw.mlir:13731:13
  wire [31:0]     _T_1694;	// matmul/matmul-hw.mlir:13730:13
  wire            _T_1695;	// matmul/matmul-hw.mlir:13729:13
  wire            _T_1696;	// matmul/matmul-hw.mlir:13728:13
  wire [31:0]     _T_1697;	// matmul/matmul-hw.mlir:13727:13
  wire            _T_1698;	// matmul/matmul-hw.mlir:13726:13
  wire            _T_1699;	// matmul/matmul-hw.mlir:13725:13
  wire [31:0]     _T_1700;	// matmul/matmul-hw.mlir:13724:13
  wire            _T_1701;	// matmul/matmul-hw.mlir:13723:13
  wire            _T_1702;	// matmul/matmul-hw.mlir:13722:13
  wire [31:0]     _T_1703;	// matmul/matmul-hw.mlir:13721:13
  wire            _T_1704;	// matmul/matmul-hw.mlir:13720:13
  wire            _T_1705;	// matmul/matmul-hw.mlir:13719:13
  wire [31:0]     _T_1706;	// matmul/matmul-hw.mlir:13718:13
  wire            _T_1707;	// matmul/matmul-hw.mlir:13717:13
  wire            _T_1708;	// matmul/matmul-hw.mlir:13716:13
  wire [31:0]     _T_1709;	// matmul/matmul-hw.mlir:13715:13
  wire            _T_1710;	// matmul/matmul-hw.mlir:13714:13
  wire            _T_1711;	// matmul/matmul-hw.mlir:13713:13
  wire [31:0]     _T_1712;	// matmul/matmul-hw.mlir:13712:13
  wire            _T_1713;	// matmul/matmul-hw.mlir:13711:13
  wire            _T_1714;	// matmul/matmul-hw.mlir:13710:13
  wire [31:0]     _T_1715;	// matmul/matmul-hw.mlir:13709:13
  wire            _T_1716;	// matmul/matmul-hw.mlir:13708:13
  wire            _T_1717;	// matmul/matmul-hw.mlir:13707:13
  wire [31:0]     _T_1718;	// matmul/matmul-hw.mlir:13706:13
  wire            _T_1719;	// matmul/matmul-hw.mlir:13705:13
  wire            _T_1720;	// matmul/matmul-hw.mlir:13704:13
  wire [31:0]     _T_1721;	// matmul/matmul-hw.mlir:13703:13
  wire            _T_1722;	// matmul/matmul-hw.mlir:13702:13
  wire            _T_1723;	// matmul/matmul-hw.mlir:13701:13
  wire [31:0]     _T_1724;	// matmul/matmul-hw.mlir:13700:13
  wire            _T_1725;	// matmul/matmul-hw.mlir:13699:13
  wire            _T_1726;	// matmul/matmul-hw.mlir:13698:13
  wire [31:0]     _T_1727;	// matmul/matmul-hw.mlir:13697:13
  wire            _T_1728;	// matmul/matmul-hw.mlir:13696:13
  wire            _T_1729;	// matmul/matmul-hw.mlir:13695:13
  wire [31:0]     _T_1730;	// matmul/matmul-hw.mlir:13679:13
  wire            _T_1731;	// matmul/matmul-hw.mlir:13678:13
  wire            _T_1732;	// matmul/matmul-hw.mlir:13677:13
  wire [31:0]     _T_1733;	// matmul/matmul-hw.mlir:13676:13
  wire            _T_1734;	// matmul/matmul-hw.mlir:13675:13
  wire            _T_1735;	// matmul/matmul-hw.mlir:13674:13
  wire [31:0]     _T_1736;	// matmul/matmul-hw.mlir:13673:13
  wire            _T_1737;	// matmul/matmul-hw.mlir:13672:13
  wire            _T_1738;	// matmul/matmul-hw.mlir:13671:13
  wire [31:0]     _T_1739;	// matmul/matmul-hw.mlir:13670:13
  wire            _T_1740;	// matmul/matmul-hw.mlir:13669:13
  wire            _T_1741;	// matmul/matmul-hw.mlir:13668:13
  wire [31:0]     _T_1742;	// matmul/matmul-hw.mlir:13667:13
  wire            _T_1743;	// matmul/matmul-hw.mlir:13666:13
  wire            _T_1744;	// matmul/matmul-hw.mlir:13665:13
  wire [31:0]     _T_1745;	// matmul/matmul-hw.mlir:13664:13
  wire            _T_1746;	// matmul/matmul-hw.mlir:13663:13
  wire            _T_1747;	// matmul/matmul-hw.mlir:13662:13
  wire [31:0]     _T_1748;	// matmul/matmul-hw.mlir:13661:13
  wire            _T_1749;	// matmul/matmul-hw.mlir:13660:13
  wire            _T_1750;	// matmul/matmul-hw.mlir:13659:13
  wire [31:0]     _T_1751;	// matmul/matmul-hw.mlir:13658:13
  wire            _T_1752;	// matmul/matmul-hw.mlir:13657:13
  wire            _T_1753;	// matmul/matmul-hw.mlir:13656:13
  wire [31:0]     _T_1754;	// matmul/matmul-hw.mlir:13655:13
  wire            _T_1755;	// matmul/matmul-hw.mlir:13654:13
  wire            _T_1756;	// matmul/matmul-hw.mlir:13653:13
  wire [31:0]     _T_1757;	// matmul/matmul-hw.mlir:13652:13
  wire            _T_1758;	// matmul/matmul-hw.mlir:13651:13
  wire            _T_1759;	// matmul/matmul-hw.mlir:13650:13
  wire [31:0]     _T_1760;	// matmul/matmul-hw.mlir:13649:13
  wire            _T_1761;	// matmul/matmul-hw.mlir:13648:13
  wire            _T_1762;	// matmul/matmul-hw.mlir:13647:13
  wire [31:0]     _T_1763;	// matmul/matmul-hw.mlir:13646:13
  wire            _T_1764;	// matmul/matmul-hw.mlir:13645:13
  wire            _T_1765;	// matmul/matmul-hw.mlir:13644:13
  wire [31:0]     _T_1766;	// matmul/matmul-hw.mlir:13643:13
  wire            _T_1767;	// matmul/matmul-hw.mlir:13642:13
  wire            _T_1768;	// matmul/matmul-hw.mlir:13641:13
  wire [31:0]     _T_1769;	// matmul/matmul-hw.mlir:13640:13
  wire            _T_1770;	// matmul/matmul-hw.mlir:13639:13
  wire            _T_1771;	// matmul/matmul-hw.mlir:13638:13
  wire [31:0]     _T_1772;	// matmul/matmul-hw.mlir:13637:13
  wire            _T_1773;	// matmul/matmul-hw.mlir:13636:13
  wire            _T_1774;	// matmul/matmul-hw.mlir:13635:12
  wire [31:0]     _T_1775;	// matmul/matmul-hw.mlir:13634:12
  wire            _T_1776;	// matmul/matmul-hw.mlir:13633:12
  wire            _T_1777;	// matmul/matmul-hw.mlir:13632:12
  wire [31:0]     _T_1778;	// matmul/matmul-hw.mlir:13616:12
  wire            _T_1779;	// matmul/matmul-hw.mlir:13615:12
  wire            _T_1780;	// matmul/matmul-hw.mlir:13614:12
  wire [31:0]     _T_1781;	// matmul/matmul-hw.mlir:13613:12
  wire            _T_1782;	// matmul/matmul-hw.mlir:13612:12
  wire            _T_1783;	// matmul/matmul-hw.mlir:13611:12
  wire [31:0]     _T_1784;	// matmul/matmul-hw.mlir:13610:12
  wire            _T_1785;	// matmul/matmul-hw.mlir:13609:12
  wire            _T_1786;	// matmul/matmul-hw.mlir:13608:12
  wire [31:0]     _T_1787;	// matmul/matmul-hw.mlir:13607:12
  wire            _T_1788;	// matmul/matmul-hw.mlir:13606:12
  wire            _T_1789;	// matmul/matmul-hw.mlir:13605:12
  wire [31:0]     _T_1790;	// matmul/matmul-hw.mlir:13604:12
  wire            _T_1791;	// matmul/matmul-hw.mlir:13603:12
  wire            _T_1792;	// matmul/matmul-hw.mlir:13602:12
  wire [31:0]     _T_1793;	// matmul/matmul-hw.mlir:13601:12
  wire            _T_1794;	// matmul/matmul-hw.mlir:13600:12
  wire            _T_1795;	// matmul/matmul-hw.mlir:13599:12
  wire [31:0]     _T_1796;	// matmul/matmul-hw.mlir:13598:12
  wire            _T_1797;	// matmul/matmul-hw.mlir:13597:12
  wire            _T_1798;	// matmul/matmul-hw.mlir:13596:12
  wire [31:0]     _T_1799;	// matmul/matmul-hw.mlir:13595:12
  wire            _T_1800;	// matmul/matmul-hw.mlir:13594:12
  wire            _T_1801;	// matmul/matmul-hw.mlir:13593:12
  wire [31:0]     _T_1802;	// matmul/matmul-hw.mlir:13592:12
  wire            _T_1803;	// matmul/matmul-hw.mlir:13591:12
  wire            _T_1804;	// matmul/matmul-hw.mlir:13590:12
  wire [31:0]     _T_1805;	// matmul/matmul-hw.mlir:13589:12
  wire            _T_1806;	// matmul/matmul-hw.mlir:13588:12
  wire            _T_1807;	// matmul/matmul-hw.mlir:13587:12
  wire [31:0]     _T_1808;	// matmul/matmul-hw.mlir:13586:12
  wire            _T_1809;	// matmul/matmul-hw.mlir:13585:12
  wire            _T_1810;	// matmul/matmul-hw.mlir:13584:12
  wire [31:0]     _T_1811;	// matmul/matmul-hw.mlir:13583:12
  wire            _T_1812;	// matmul/matmul-hw.mlir:13582:12
  wire            _T_1813;	// matmul/matmul-hw.mlir:13581:12
  wire [31:0]     _T_1814;	// matmul/matmul-hw.mlir:13580:12
  wire            _T_1815;	// matmul/matmul-hw.mlir:13579:12
  wire            _T_1816;	// matmul/matmul-hw.mlir:13578:12
  wire [31:0]     _T_1817;	// matmul/matmul-hw.mlir:13577:12
  wire            _T_1818;	// matmul/matmul-hw.mlir:13576:12
  wire            _T_1819;	// matmul/matmul-hw.mlir:13575:12
  wire [31:0]     _T_1820;	// matmul/matmul-hw.mlir:13574:12
  wire            _T_1821;	// matmul/matmul-hw.mlir:13573:12
  wire            _T_1822;	// matmul/matmul-hw.mlir:13572:12
  wire [31:0]     _T_1823;	// matmul/matmul-hw.mlir:13571:12
  wire            _T_1824;	// matmul/matmul-hw.mlir:13570:12
  wire            _T_1825;	// matmul/matmul-hw.mlir:13569:12
  wire [31:0]     _T_1826;	// matmul/matmul-hw.mlir:13553:12
  wire            _T_1827;	// matmul/matmul-hw.mlir:13552:12
  wire            _T_1828;	// matmul/matmul-hw.mlir:13551:12
  wire [31:0]     _T_1829;	// matmul/matmul-hw.mlir:13550:12
  wire            _T_1830;	// matmul/matmul-hw.mlir:13549:12
  wire            _T_1831;	// matmul/matmul-hw.mlir:13548:12
  wire [31:0]     _T_1832;	// matmul/matmul-hw.mlir:13547:12
  wire            _T_1833;	// matmul/matmul-hw.mlir:13546:12
  wire            _T_1834;	// matmul/matmul-hw.mlir:13545:12
  wire [31:0]     _T_1835;	// matmul/matmul-hw.mlir:13544:12
  wire            _T_1836;	// matmul/matmul-hw.mlir:13543:12
  wire            _T_1837;	// matmul/matmul-hw.mlir:13542:12
  wire [31:0]     _T_1838;	// matmul/matmul-hw.mlir:13541:12
  wire            _T_1839;	// matmul/matmul-hw.mlir:13540:12
  wire            _T_1840;	// matmul/matmul-hw.mlir:13539:12
  wire [31:0]     _T_1841;	// matmul/matmul-hw.mlir:13538:12
  wire            _T_1842;	// matmul/matmul-hw.mlir:13537:12
  wire            _T_1843;	// matmul/matmul-hw.mlir:13536:12
  wire [31:0]     _T_1844;	// matmul/matmul-hw.mlir:13535:12
  wire            _T_1845;	// matmul/matmul-hw.mlir:13534:12
  wire            _T_1846;	// matmul/matmul-hw.mlir:13533:12
  wire [31:0]     _T_1847;	// matmul/matmul-hw.mlir:13532:12
  wire            _T_1848;	// matmul/matmul-hw.mlir:13531:12
  wire            _T_1849;	// matmul/matmul-hw.mlir:13530:12
  wire [31:0]     _T_1850;	// matmul/matmul-hw.mlir:13529:12
  wire            _T_1851;	// matmul/matmul-hw.mlir:13528:12
  wire            _T_1852;	// matmul/matmul-hw.mlir:13527:12
  wire [31:0]     _T_1853;	// matmul/matmul-hw.mlir:13526:12
  wire            _T_1854;	// matmul/matmul-hw.mlir:13525:12
  wire            _T_1855;	// matmul/matmul-hw.mlir:13524:12
  wire [31:0]     _T_1856;	// matmul/matmul-hw.mlir:13523:12
  wire            _T_1857;	// matmul/matmul-hw.mlir:13522:12
  wire            _T_1858;	// matmul/matmul-hw.mlir:13521:12
  wire [31:0]     _T_1859;	// matmul/matmul-hw.mlir:13520:12
  wire            _T_1860;	// matmul/matmul-hw.mlir:13519:12
  wire            _T_1861;	// matmul/matmul-hw.mlir:13518:12
  wire [31:0]     _T_1862;	// matmul/matmul-hw.mlir:13517:12
  wire            _T_1863;	// matmul/matmul-hw.mlir:13516:12
  wire            _T_1864;	// matmul/matmul-hw.mlir:13515:12
  wire [31:0]     _T_1865;	// matmul/matmul-hw.mlir:13514:12
  wire            _T_1866;	// matmul/matmul-hw.mlir:13513:12
  wire            _T_1867;	// matmul/matmul-hw.mlir:13512:12
  wire [31:0]     _T_1868;	// matmul/matmul-hw.mlir:13511:12
  wire            _T_1869;	// matmul/matmul-hw.mlir:13510:12
  wire            _T_1870;	// matmul/matmul-hw.mlir:13509:12
  wire [31:0]     _T_1871;	// matmul/matmul-hw.mlir:13508:12
  wire            _T_1872;	// matmul/matmul-hw.mlir:13507:12
  wire            _T_1873;	// matmul/matmul-hw.mlir:13506:12
  wire [31:0]     _T_1874;	// matmul/matmul-hw.mlir:13490:12
  wire            _T_1875;	// matmul/matmul-hw.mlir:13489:12
  wire            _T_1876;	// matmul/matmul-hw.mlir:13488:12
  wire [31:0]     _T_1877;	// matmul/matmul-hw.mlir:13487:12
  wire            _T_1878;	// matmul/matmul-hw.mlir:13486:12
  wire            _T_1879;	// matmul/matmul-hw.mlir:13485:12
  wire [31:0]     _T_1880;	// matmul/matmul-hw.mlir:13484:12
  wire            _T_1881;	// matmul/matmul-hw.mlir:13483:12
  wire            _T_1882;	// matmul/matmul-hw.mlir:13482:12
  wire [31:0]     _T_1883;	// matmul/matmul-hw.mlir:13481:12
  wire            _T_1884;	// matmul/matmul-hw.mlir:13480:12
  wire            _T_1885;	// matmul/matmul-hw.mlir:13479:12
  wire [31:0]     _T_1886;	// matmul/matmul-hw.mlir:13478:12
  wire            _T_1887;	// matmul/matmul-hw.mlir:13477:12
  wire            _T_1888;	// matmul/matmul-hw.mlir:13476:12
  wire [31:0]     _T_1889;	// matmul/matmul-hw.mlir:13475:12
  wire            _T_1890;	// matmul/matmul-hw.mlir:13474:12
  wire            _T_1891;	// matmul/matmul-hw.mlir:13473:12
  wire [31:0]     _T_1892;	// matmul/matmul-hw.mlir:13472:12
  wire            _T_1893;	// matmul/matmul-hw.mlir:13471:12
  wire            _T_1894;	// matmul/matmul-hw.mlir:13470:12
  wire [31:0]     _T_1895;	// matmul/matmul-hw.mlir:13469:12
  wire            _T_1896;	// matmul/matmul-hw.mlir:13468:12
  wire            _T_1897;	// matmul/matmul-hw.mlir:13467:12
  wire [31:0]     _T_1898;	// matmul/matmul-hw.mlir:13466:12
  wire            _T_1899;	// matmul/matmul-hw.mlir:13465:12
  wire            _T_1900;	// matmul/matmul-hw.mlir:13464:12
  wire [31:0]     _T_1901;	// matmul/matmul-hw.mlir:13463:12
  wire            _T_1902;	// matmul/matmul-hw.mlir:13462:12
  wire            _T_1903;	// matmul/matmul-hw.mlir:13461:12
  wire [31:0]     _T_1904;	// matmul/matmul-hw.mlir:13460:12
  wire            _T_1905;	// matmul/matmul-hw.mlir:13459:12
  wire            _T_1906;	// matmul/matmul-hw.mlir:13458:12
  wire [31:0]     _T_1907;	// matmul/matmul-hw.mlir:13457:12
  wire            _T_1908;	// matmul/matmul-hw.mlir:13456:12
  wire            _T_1909;	// matmul/matmul-hw.mlir:13455:12
  wire [31:0]     _T_1910;	// matmul/matmul-hw.mlir:13454:12
  wire            _T_1911;	// matmul/matmul-hw.mlir:13453:12
  wire            _T_1912;	// matmul/matmul-hw.mlir:13452:12
  wire [31:0]     _T_1913;	// matmul/matmul-hw.mlir:13451:12
  wire            _T_1914;	// matmul/matmul-hw.mlir:13450:12
  wire            _T_1915;	// matmul/matmul-hw.mlir:13449:12
  wire [31:0]     _T_1916;	// matmul/matmul-hw.mlir:13448:12
  wire            _T_1917;	// matmul/matmul-hw.mlir:13447:12
  wire            _T_1918;	// matmul/matmul-hw.mlir:13446:12
  wire [31:0]     _T_1919;	// matmul/matmul-hw.mlir:13445:12
  wire            _T_1920;	// matmul/matmul-hw.mlir:13444:12
  wire            _T_1921;	// matmul/matmul-hw.mlir:13443:12
  wire [31:0]     _T_1922;	// matmul/matmul-hw.mlir:13427:12
  wire            _T_1923;	// matmul/matmul-hw.mlir:13426:12
  wire            _T_1924;	// matmul/matmul-hw.mlir:13425:12
  wire [31:0]     _T_1925;	// matmul/matmul-hw.mlir:13424:12
  wire            _T_1926;	// matmul/matmul-hw.mlir:13423:12
  wire            _T_1927;	// matmul/matmul-hw.mlir:13422:12
  wire [31:0]     _T_1928;	// matmul/matmul-hw.mlir:13421:12
  wire            _T_1929;	// matmul/matmul-hw.mlir:13420:12
  wire            _T_1930;	// matmul/matmul-hw.mlir:13419:12
  wire [31:0]     _T_1931;	// matmul/matmul-hw.mlir:13418:12
  wire            _T_1932;	// matmul/matmul-hw.mlir:13417:12
  wire            _T_1933;	// matmul/matmul-hw.mlir:13416:12
  wire [31:0]     _T_1934;	// matmul/matmul-hw.mlir:13415:12
  wire            _T_1935;	// matmul/matmul-hw.mlir:13414:12
  wire            _T_1936;	// matmul/matmul-hw.mlir:13413:12
  wire [31:0]     _T_1937;	// matmul/matmul-hw.mlir:13412:12
  wire            _T_1938;	// matmul/matmul-hw.mlir:13411:12
  wire            _T_1939;	// matmul/matmul-hw.mlir:13410:12
  wire [31:0]     _T_1940;	// matmul/matmul-hw.mlir:13409:12
  wire            _T_1941;	// matmul/matmul-hw.mlir:13408:12
  wire            _T_1942;	// matmul/matmul-hw.mlir:13407:12
  wire [31:0]     _T_1943;	// matmul/matmul-hw.mlir:13406:12
  wire            _T_1944;	// matmul/matmul-hw.mlir:13405:12
  wire            _T_1945;	// matmul/matmul-hw.mlir:13404:12
  wire [31:0]     _T_1946;	// matmul/matmul-hw.mlir:13403:12
  wire            _T_1947;	// matmul/matmul-hw.mlir:13402:12
  wire            _T_1948;	// matmul/matmul-hw.mlir:13401:12
  wire [31:0]     _T_1949;	// matmul/matmul-hw.mlir:13400:12
  wire            _T_1950;	// matmul/matmul-hw.mlir:13399:12
  wire            _T_1951;	// matmul/matmul-hw.mlir:13398:12
  wire [31:0]     _T_1952;	// matmul/matmul-hw.mlir:13397:12
  wire            _T_1953;	// matmul/matmul-hw.mlir:13396:12
  wire            _T_1954;	// matmul/matmul-hw.mlir:13395:12
  wire [31:0]     _T_1955;	// matmul/matmul-hw.mlir:13394:12
  wire            _T_1956;	// matmul/matmul-hw.mlir:13393:12
  wire            _T_1957;	// matmul/matmul-hw.mlir:13392:12
  wire [31:0]     _T_1958;	// matmul/matmul-hw.mlir:13391:12
  wire            _T_1959;	// matmul/matmul-hw.mlir:13390:12
  wire            _T_1960;	// matmul/matmul-hw.mlir:13389:12
  wire [31:0]     _T_1961;	// matmul/matmul-hw.mlir:13388:12
  wire            _T_1962;	// matmul/matmul-hw.mlir:13387:12
  wire            _T_1963;	// matmul/matmul-hw.mlir:13386:12
  wire [31:0]     _T_1964;	// matmul/matmul-hw.mlir:13385:12
  wire            _T_1965;	// matmul/matmul-hw.mlir:13384:12
  wire            _T_1966;	// matmul/matmul-hw.mlir:13383:12
  wire [31:0]     _T_1967;	// matmul/matmul-hw.mlir:13382:12
  wire            _T_1968;	// matmul/matmul-hw.mlir:13381:12
  wire            _T_1969;	// matmul/matmul-hw.mlir:13380:12
  wire [31:0]     _T_1970;	// matmul/matmul-hw.mlir:13364:12
  wire            _T_1971;	// matmul/matmul-hw.mlir:13363:12
  wire            _T_1972;	// matmul/matmul-hw.mlir:13362:12
  wire [31:0]     _T_1973;	// matmul/matmul-hw.mlir:13361:12
  wire            _T_1974;	// matmul/matmul-hw.mlir:13360:12
  wire            _T_1975;	// matmul/matmul-hw.mlir:13359:12
  wire [31:0]     _T_1976;	// matmul/matmul-hw.mlir:13358:12
  wire            _T_1977;	// matmul/matmul-hw.mlir:13357:12
  wire            _T_1978;	// matmul/matmul-hw.mlir:13356:12
  wire [31:0]     _T_1979;	// matmul/matmul-hw.mlir:13355:12
  wire            _T_1980;	// matmul/matmul-hw.mlir:13354:12
  wire            _T_1981;	// matmul/matmul-hw.mlir:13353:12
  wire [31:0]     _T_1982;	// matmul/matmul-hw.mlir:13352:12
  wire            _T_1983;	// matmul/matmul-hw.mlir:13351:12
  wire            _T_1984;	// matmul/matmul-hw.mlir:13350:12
  wire [31:0]     _T_1985;	// matmul/matmul-hw.mlir:13349:12
  wire            _T_1986;	// matmul/matmul-hw.mlir:13348:12
  wire            _T_1987;	// matmul/matmul-hw.mlir:13347:12
  wire [31:0]     _T_1988;	// matmul/matmul-hw.mlir:13346:12
  wire            _T_1989;	// matmul/matmul-hw.mlir:13345:12
  wire            _T_1990;	// matmul/matmul-hw.mlir:13344:12
  wire [31:0]     _T_1991;	// matmul/matmul-hw.mlir:13343:12
  wire            _T_1992;	// matmul/matmul-hw.mlir:13342:12
  wire            _T_1993;	// matmul/matmul-hw.mlir:13341:12
  wire [31:0]     _T_1994;	// matmul/matmul-hw.mlir:13340:12
  wire            _T_1995;	// matmul/matmul-hw.mlir:13339:12
  wire            _T_1996;	// matmul/matmul-hw.mlir:13338:12
  wire [31:0]     _T_1997;	// matmul/matmul-hw.mlir:13337:12
  wire            _T_1998;	// matmul/matmul-hw.mlir:13336:12
  wire            _T_1999;	// matmul/matmul-hw.mlir:13335:12
  wire [31:0]     _T_2000;	// matmul/matmul-hw.mlir:13334:12
  wire            _T_2001;	// matmul/matmul-hw.mlir:13333:12
  wire            _T_2002;	// matmul/matmul-hw.mlir:13332:12
  wire [31:0]     _T_2003;	// matmul/matmul-hw.mlir:13331:12
  wire            _T_2004;	// matmul/matmul-hw.mlir:13330:12
  wire            _T_2005;	// matmul/matmul-hw.mlir:13329:12
  wire [31:0]     _T_2006;	// matmul/matmul-hw.mlir:13328:12
  wire            _T_2007;	// matmul/matmul-hw.mlir:13327:12
  wire            _T_2008;	// matmul/matmul-hw.mlir:13326:12
  wire [31:0]     _T_2009;	// matmul/matmul-hw.mlir:13325:12
  wire            _T_2010;	// matmul/matmul-hw.mlir:13324:12
  wire            _T_2011;	// matmul/matmul-hw.mlir:13323:12
  wire [31:0]     _T_2012;	// matmul/matmul-hw.mlir:13322:12
  wire            _T_2013;	// matmul/matmul-hw.mlir:13321:12
  wire            _T_2014;	// matmul/matmul-hw.mlir:13320:12
  wire [31:0]     _T_2015;	// matmul/matmul-hw.mlir:13319:12
  wire            _T_2016;	// matmul/matmul-hw.mlir:13318:12
  wire            _T_2017;	// matmul/matmul-hw.mlir:13317:12
  wire [31:0]     _T_2018;	// matmul/matmul-hw.mlir:13301:12
  wire            _T_2019;	// matmul/matmul-hw.mlir:13300:12
  wire            _T_2020;	// matmul/matmul-hw.mlir:13299:12
  wire [31:0]     _T_2021;	// matmul/matmul-hw.mlir:13298:12
  wire            _T_2022;	// matmul/matmul-hw.mlir:13297:12
  wire            _T_2023;	// matmul/matmul-hw.mlir:13296:12
  wire [31:0]     _T_2024;	// matmul/matmul-hw.mlir:13295:12
  wire            _T_2025;	// matmul/matmul-hw.mlir:13294:12
  wire            _T_2026;	// matmul/matmul-hw.mlir:13293:12
  wire [31:0]     _T_2027;	// matmul/matmul-hw.mlir:13292:12
  wire            _T_2028;	// matmul/matmul-hw.mlir:13291:12
  wire            _T_2029;	// matmul/matmul-hw.mlir:13290:12
  wire [31:0]     _T_2030;	// matmul/matmul-hw.mlir:13289:12
  wire            _T_2031;	// matmul/matmul-hw.mlir:13288:12
  wire            _T_2032;	// matmul/matmul-hw.mlir:13287:12
  wire [31:0]     _T_2033;	// matmul/matmul-hw.mlir:13286:12
  wire            _T_2034;	// matmul/matmul-hw.mlir:13285:12
  wire            _T_2035;	// matmul/matmul-hw.mlir:13284:12
  wire [31:0]     _T_2036;	// matmul/matmul-hw.mlir:13283:12
  wire            _T_2037;	// matmul/matmul-hw.mlir:13282:12
  wire            _T_2038;	// matmul/matmul-hw.mlir:13281:12
  wire [31:0]     _T_2039;	// matmul/matmul-hw.mlir:13280:12
  wire            _T_2040;	// matmul/matmul-hw.mlir:13279:12
  wire            _T_2041;	// matmul/matmul-hw.mlir:13278:12
  wire [31:0]     _T_2042;	// matmul/matmul-hw.mlir:13277:12
  wire            _T_2043;	// matmul/matmul-hw.mlir:13276:12
  wire            _T_2044;	// matmul/matmul-hw.mlir:13275:12
  wire [31:0]     _T_2045;	// matmul/matmul-hw.mlir:13274:12
  wire            _T_2046;	// matmul/matmul-hw.mlir:13273:12
  wire            _T_2047;	// matmul/matmul-hw.mlir:13272:12
  wire [31:0]     _T_2048;	// matmul/matmul-hw.mlir:13271:12
  wire            _T_2049;	// matmul/matmul-hw.mlir:13270:12
  wire            _T_2050;	// matmul/matmul-hw.mlir:13269:12
  wire [31:0]     _T_2051;	// matmul/matmul-hw.mlir:13268:12
  wire            _T_2052;	// matmul/matmul-hw.mlir:13267:12
  wire            _T_2053;	// matmul/matmul-hw.mlir:13266:12
  wire [31:0]     _T_2054;	// matmul/matmul-hw.mlir:13265:12
  wire            _T_2055;	// matmul/matmul-hw.mlir:13264:12
  wire            _T_2056;	// matmul/matmul-hw.mlir:13263:12
  wire [31:0]     _T_2057;	// matmul/matmul-hw.mlir:13262:12
  wire            _T_2058;	// matmul/matmul-hw.mlir:13261:12
  wire            _T_2059;	// matmul/matmul-hw.mlir:13260:12
  wire [31:0]     _T_2060;	// matmul/matmul-hw.mlir:13259:12
  wire            _T_2061;	// matmul/matmul-hw.mlir:13258:12
  wire            _T_2062;	// matmul/matmul-hw.mlir:13257:12
  wire [31:0]     _T_2063;	// matmul/matmul-hw.mlir:13256:12
  wire            _T_2064;	// matmul/matmul-hw.mlir:13255:12
  wire            _T_2065;	// matmul/matmul-hw.mlir:13254:12
  wire [31:0]     _T_2066;	// matmul/matmul-hw.mlir:13238:12
  wire            _T_2067;	// matmul/matmul-hw.mlir:13237:12
  wire            _T_2068;	// matmul/matmul-hw.mlir:13236:12
  wire [31:0]     _T_2069;	// matmul/matmul-hw.mlir:13235:12
  wire            _T_2070;	// matmul/matmul-hw.mlir:13234:12
  wire            _T_2071;	// matmul/matmul-hw.mlir:13233:12
  wire [31:0]     _T_2072;	// matmul/matmul-hw.mlir:13232:12
  wire            _T_2073;	// matmul/matmul-hw.mlir:13231:12
  wire            _T_2074;	// matmul/matmul-hw.mlir:13230:12
  wire [31:0]     _T_2075;	// matmul/matmul-hw.mlir:13229:12
  wire            _T_2076;	// matmul/matmul-hw.mlir:13228:12
  wire            _T_2077;	// matmul/matmul-hw.mlir:13227:12
  wire [31:0]     _T_2078;	// matmul/matmul-hw.mlir:13226:12
  wire            _T_2079;	// matmul/matmul-hw.mlir:13225:12
  wire            _T_2080;	// matmul/matmul-hw.mlir:13224:12
  wire [31:0]     _T_2081;	// matmul/matmul-hw.mlir:13223:12
  wire            _T_2082;	// matmul/matmul-hw.mlir:13222:12
  wire            _T_2083;	// matmul/matmul-hw.mlir:13221:12
  wire [31:0]     _T_2084;	// matmul/matmul-hw.mlir:13220:12
  wire            _T_2085;	// matmul/matmul-hw.mlir:13219:12
  wire            _T_2086;	// matmul/matmul-hw.mlir:13218:12
  wire [31:0]     _T_2087;	// matmul/matmul-hw.mlir:13217:12
  wire            _T_2088;	// matmul/matmul-hw.mlir:13216:12
  wire            _T_2089;	// matmul/matmul-hw.mlir:13215:12
  wire [31:0]     _T_2090;	// matmul/matmul-hw.mlir:13214:12
  wire            _T_2091;	// matmul/matmul-hw.mlir:13213:12
  wire            _T_2092;	// matmul/matmul-hw.mlir:13212:12
  wire [31:0]     _T_2093;	// matmul/matmul-hw.mlir:13211:12
  wire            _T_2094;	// matmul/matmul-hw.mlir:13210:12
  wire            _T_2095;	// matmul/matmul-hw.mlir:13209:12
  wire [31:0]     _T_2096;	// matmul/matmul-hw.mlir:13208:12
  wire            _T_2097;	// matmul/matmul-hw.mlir:13207:12
  wire            _T_2098;	// matmul/matmul-hw.mlir:13206:12
  wire [31:0]     _T_2099;	// matmul/matmul-hw.mlir:13205:12
  wire            _T_2100;	// matmul/matmul-hw.mlir:13204:12
  wire            _T_2101;	// matmul/matmul-hw.mlir:13203:12
  wire [31:0]     _T_2102;	// matmul/matmul-hw.mlir:13202:12
  wire            _T_2103;	// matmul/matmul-hw.mlir:13201:12
  wire            _T_2104;	// matmul/matmul-hw.mlir:13200:12
  wire [31:0]     _T_2105;	// matmul/matmul-hw.mlir:13199:12
  wire            _T_2106;	// matmul/matmul-hw.mlir:13198:12
  wire            _T_2107;	// matmul/matmul-hw.mlir:13197:12
  wire [31:0]     _T_2108;	// matmul/matmul-hw.mlir:13196:12
  wire            _T_2109;	// matmul/matmul-hw.mlir:13195:12
  wire            _T_2110;	// matmul/matmul-hw.mlir:13194:12
  wire [31:0]     _T_2111;	// matmul/matmul-hw.mlir:13182:12
  wire            _T_2112;	// matmul/matmul-hw.mlir:13181:12
  wire            _T_2113;	// matmul/matmul-hw.mlir:13150:12
  wire [3:0]      _T_2114;	// matmul/matmul-hw.mlir:13149:12
  wire            _T_2115;	// matmul/matmul-hw.mlir:13148:12
  wire [31:0]     _T_2116;	// matmul/matmul-hw.mlir:13136:12
  wire            _T_2117;	// matmul/matmul-hw.mlir:13135:12
  wire            _T_2118;	// matmul/matmul-hw.mlir:13104:12
  wire [3:0]      _T_2119;	// matmul/matmul-hw.mlir:13103:12
  wire            _T_2120;	// matmul/matmul-hw.mlir:13102:12
  wire [31:0]     _T_2121;	// matmul/matmul-hw.mlir:13090:12
  wire            _T_2122;	// matmul/matmul-hw.mlir:13089:12
  wire            _T_2123;	// matmul/matmul-hw.mlir:13058:12
  wire [3:0]      _T_2124;	// matmul/matmul-hw.mlir:13057:12
  wire            _T_2125;	// matmul/matmul-hw.mlir:13056:12
  wire [31:0]     _T_2126;	// matmul/matmul-hw.mlir:13044:12
  wire            _T_2127;	// matmul/matmul-hw.mlir:13043:12
  wire            _T_2128;	// matmul/matmul-hw.mlir:13012:12
  wire [3:0]      _T_2129;	// matmul/matmul-hw.mlir:13011:12
  wire            _T_2130;	// matmul/matmul-hw.mlir:13010:12
  wire [31:0]     _T_2131;	// matmul/matmul-hw.mlir:12998:12
  wire            _T_2132;	// matmul/matmul-hw.mlir:12997:12
  wire            _T_2133;	// matmul/matmul-hw.mlir:12966:12
  wire [3:0]      _T_2134;	// matmul/matmul-hw.mlir:12965:12
  wire            _T_2135;	// matmul/matmul-hw.mlir:12964:12
  wire [31:0]     _T_2136;	// matmul/matmul-hw.mlir:12952:12
  wire            _T_2137;	// matmul/matmul-hw.mlir:12951:12
  wire            _T_2138;	// matmul/matmul-hw.mlir:12920:12
  wire [3:0]      _T_2139;	// matmul/matmul-hw.mlir:12919:12
  wire            _T_2140;	// matmul/matmul-hw.mlir:12918:12
  wire [31:0]     _T_2141;	// matmul/matmul-hw.mlir:12906:12
  wire            _T_2142;	// matmul/matmul-hw.mlir:12905:12
  wire            _T_2143;	// matmul/matmul-hw.mlir:12874:12
  wire [3:0]      _T_2144;	// matmul/matmul-hw.mlir:12873:12
  wire            _T_2145;	// matmul/matmul-hw.mlir:12872:12
  wire [31:0]     _T_2146;	// matmul/matmul-hw.mlir:12860:12
  wire            _T_2147;	// matmul/matmul-hw.mlir:12859:12
  wire            _T_2148;	// matmul/matmul-hw.mlir:12828:12
  wire [3:0]      _T_2149;	// matmul/matmul-hw.mlir:12827:12
  wire            _T_2150;	// matmul/matmul-hw.mlir:12826:12
  wire [31:0]     _T_2151;	// matmul/matmul-hw.mlir:12814:12
  wire            _T_2152;	// matmul/matmul-hw.mlir:12813:12
  wire            _T_2153;	// matmul/matmul-hw.mlir:12782:12
  wire [3:0]      _T_2154;	// matmul/matmul-hw.mlir:12781:12
  wire            _T_2155;	// matmul/matmul-hw.mlir:12780:12
  wire [31:0]     _T_2156;	// matmul/matmul-hw.mlir:12768:12
  wire            _T_2157;	// matmul/matmul-hw.mlir:12767:12
  wire            _T_2158;	// matmul/matmul-hw.mlir:12736:12
  wire [3:0]      _T_2159;	// matmul/matmul-hw.mlir:12735:12
  wire            _T_2160;	// matmul/matmul-hw.mlir:12734:12
  wire [31:0]     _T_2161;	// matmul/matmul-hw.mlir:12722:12
  wire            _T_2162;	// matmul/matmul-hw.mlir:12721:12
  wire            _T_2163;	// matmul/matmul-hw.mlir:12690:12
  wire [3:0]      _T_2164;	// matmul/matmul-hw.mlir:12689:12
  wire            _T_2165;	// matmul/matmul-hw.mlir:12688:12
  wire [31:0]     _T_2166;	// matmul/matmul-hw.mlir:12676:12
  wire            _T_2167;	// matmul/matmul-hw.mlir:12675:12
  wire            _T_2168;	// matmul/matmul-hw.mlir:12644:12
  wire [3:0]      _T_2169;	// matmul/matmul-hw.mlir:12643:12
  wire            _T_2170;	// matmul/matmul-hw.mlir:12642:12
  wire [31:0]     _T_2171;	// matmul/matmul-hw.mlir:12630:12
  wire            _T_2172;	// matmul/matmul-hw.mlir:12629:12
  wire            _T_2173;	// matmul/matmul-hw.mlir:12598:12
  wire [3:0]      _T_2174;	// matmul/matmul-hw.mlir:12597:12
  wire            _T_2175;	// matmul/matmul-hw.mlir:12596:12
  wire [31:0]     _T_2176;	// matmul/matmul-hw.mlir:12584:12
  wire            _T_2177;	// matmul/matmul-hw.mlir:12583:12
  wire            _T_2178;	// matmul/matmul-hw.mlir:12552:12
  wire [3:0]      _T_2179;	// matmul/matmul-hw.mlir:12551:12
  wire            _T_2180;	// matmul/matmul-hw.mlir:12550:12
  wire [31:0]     _T_2181;	// matmul/matmul-hw.mlir:12538:12
  wire            _T_2182;	// matmul/matmul-hw.mlir:12537:12
  wire            _T_2183;	// matmul/matmul-hw.mlir:12506:12
  wire [3:0]      _T_2184;	// matmul/matmul-hw.mlir:12505:12
  wire            _T_2185;	// matmul/matmul-hw.mlir:12504:12
  wire [31:0]     _T_2186;	// matmul/matmul-hw.mlir:12492:12
  wire            _T_2187;	// matmul/matmul-hw.mlir:12491:12
  wire            _T_2188;	// matmul/matmul-hw.mlir:12484:12
  reg             _T_2189;	// matmul/matmul-hw.mlir:12483:12
  wire            _T_2190;	// matmul/matmul-hw.mlir:12474:12
  wire [3:0]      _T_2191;	// matmul/matmul-hw.mlir:12473:12
  wire            _T_2192;	// matmul/matmul-hw.mlir:12472:12
  wire            _T_2193;	// matmul/matmul-hw.mlir:11181:12
  wire            _T_2194;	// matmul/matmul-hw.mlir:11180:12
  wire            _T_2195;	// matmul/matmul-hw.mlir:11179:12
  wire [5:0]      _T_2196;	// matmul/matmul-hw.mlir:11172:12
  wire            _T_2197;	// matmul/matmul-hw.mlir:11171:12
  wire            _T_2198;	// matmul/matmul-hw.mlir:11168:12
  wire [31:0]     mult_inst255_result;	// matmul/matmul-hw.mlir:23520:28
  wire [31:0]     mult_inst254_result;	// matmul/matmul-hw.mlir:23490:28
  wire [31:0]     mult_inst253_result;	// matmul/matmul-hw.mlir:23460:28
  wire [31:0]     mult_inst252_result;	// matmul/matmul-hw.mlir:23430:28
  wire [31:0]     mult_inst251_result;	// matmul/matmul-hw.mlir:23400:28
  wire [31:0]     mult_inst250_result;	// matmul/matmul-hw.mlir:23370:28
  wire [31:0]     mult_inst249_result;	// matmul/matmul-hw.mlir:23340:28
  wire [31:0]     mult_inst248_result;	// matmul/matmul-hw.mlir:23310:28
  wire [31:0]     mult_inst247_result;	// matmul/matmul-hw.mlir:23280:28
  wire [31:0]     mult_inst246_result;	// matmul/matmul-hw.mlir:23250:28
  wire [31:0]     mult_inst245_result;	// matmul/matmul-hw.mlir:23220:28
  wire [31:0]     mult_inst244_result;	// matmul/matmul-hw.mlir:23190:28
  wire [31:0]     mult_inst243_result;	// matmul/matmul-hw.mlir:23160:28
  wire [31:0]     mult_inst242_result;	// matmul/matmul-hw.mlir:23130:28
  wire [31:0]     mult_inst241_result;	// matmul/matmul-hw.mlir:23100:28
  wire [31:0]     mult_inst240_result;	// matmul/matmul-hw.mlir:23070:28
  wire [31:0]     C_reg_bank16_p0_rd_data;	// matmul/matmul-hw.mlir:23065:37
  wire [31:0]     C_reg_bank15_p0_rd_data;	// matmul/matmul-hw.mlir:23064:37
  wire [31:0]     C_reg_bank14_p0_rd_data;	// matmul/matmul-hw.mlir:23063:37
  wire [31:0]     C_reg_bank13_p0_rd_data;	// matmul/matmul-hw.mlir:23062:37
  wire [31:0]     C_reg_bank12_p0_rd_data;	// matmul/matmul-hw.mlir:23061:37
  wire [31:0]     C_reg_bank11_p0_rd_data;	// matmul/matmul-hw.mlir:23060:37
  wire [31:0]     C_reg_bank10_p0_rd_data;	// matmul/matmul-hw.mlir:23059:37
  wire [31:0]     C_reg_bank9_p0_rd_data;	// matmul/matmul-hw.mlir:23058:36
  wire [31:0]     C_reg_bank8_p0_rd_data;	// matmul/matmul-hw.mlir:23057:36
  wire [31:0]     C_reg_bank7_p0_rd_data;	// matmul/matmul-hw.mlir:23056:36
  wire [31:0]     C_reg_bank6_p0_rd_data;	// matmul/matmul-hw.mlir:23055:36
  wire [31:0]     C_reg_bank5_p0_rd_data;	// matmul/matmul-hw.mlir:23054:36
  wire [31:0]     C_reg_bank4_p0_rd_data;	// matmul/matmul-hw.mlir:23053:36
  wire [31:0]     C_reg_bank3_p0_rd_data;	// matmul/matmul-hw.mlir:23052:36
  wire [31:0]     C_reg_bank2_p0_rd_data;	// matmul/matmul-hw.mlir:23051:36
  wire [31:0]     C_reg_bank1_p0_rd_data;	// matmul/matmul-hw.mlir:23050:36
  wire [31:0]     C_reg_bank0_p0_rd_data;	// matmul/matmul-hw.mlir:23049:36
  wire [31:0]     mult_inst239_result;	// matmul/matmul-hw.mlir:22910:28
  wire [31:0]     mult_inst238_result;	// matmul/matmul-hw.mlir:22880:28
  wire [31:0]     mult_inst237_result;	// matmul/matmul-hw.mlir:22850:28
  wire [31:0]     mult_inst236_result;	// matmul/matmul-hw.mlir:22820:28
  wire [31:0]     mult_inst235_result;	// matmul/matmul-hw.mlir:22790:28
  wire [31:0]     mult_inst234_result;	// matmul/matmul-hw.mlir:22760:28
  wire [31:0]     mult_inst233_result;	// matmul/matmul-hw.mlir:22730:28
  wire [31:0]     mult_inst232_result;	// matmul/matmul-hw.mlir:22700:28
  wire [31:0]     mult_inst231_result;	// matmul/matmul-hw.mlir:22670:28
  wire [31:0]     mult_inst230_result;	// matmul/matmul-hw.mlir:22640:28
  wire [31:0]     mult_inst229_result;	// matmul/matmul-hw.mlir:22610:28
  wire [31:0]     mult_inst228_result;	// matmul/matmul-hw.mlir:22580:28
  wire [31:0]     mult_inst227_result;	// matmul/matmul-hw.mlir:22550:28
  wire [31:0]     mult_inst226_result;	// matmul/matmul-hw.mlir:22520:28
  wire [31:0]     mult_inst225_result;	// matmul/matmul-hw.mlir:22490:28
  wire [31:0]     mult_inst224_result;	// matmul/matmul-hw.mlir:22460:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2199;	// matmul/matmul-hw.mlir:22455:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2200;	// matmul/matmul-hw.mlir:22454:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2201;	// matmul/matmul-hw.mlir:22453:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2202;	// matmul/matmul-hw.mlir:22452:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2203;	// matmul/matmul-hw.mlir:22451:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2204;	// matmul/matmul-hw.mlir:22450:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2205;	// matmul/matmul-hw.mlir:22449:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2206;	// matmul/matmul-hw.mlir:22448:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2207;	// matmul/matmul-hw.mlir:22447:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2208;	// matmul/matmul-hw.mlir:22446:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2209;	// matmul/matmul-hw.mlir:22445:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2210;	// matmul/matmul-hw.mlir:22444:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2211;	// matmul/matmul-hw.mlir:22443:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2212;	// matmul/matmul-hw.mlir:22442:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2213;	// matmul/matmul-hw.mlir:22441:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2214;	// matmul/matmul-hw.mlir:22440:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2215;	// matmul/matmul-hw.mlir:22439:36
  wire [31:0]     mult_inst223_result;	// matmul/matmul-hw.mlir:22300:28
  wire [31:0]     mult_inst222_result;	// matmul/matmul-hw.mlir:22270:28
  wire [31:0]     mult_inst221_result;	// matmul/matmul-hw.mlir:22240:28
  wire [31:0]     mult_inst220_result;	// matmul/matmul-hw.mlir:22210:28
  wire [31:0]     mult_inst219_result;	// matmul/matmul-hw.mlir:22180:28
  wire [31:0]     mult_inst218_result;	// matmul/matmul-hw.mlir:22150:28
  wire [31:0]     mult_inst217_result;	// matmul/matmul-hw.mlir:22120:28
  wire [31:0]     mult_inst216_result;	// matmul/matmul-hw.mlir:22090:28
  wire [31:0]     mult_inst215_result;	// matmul/matmul-hw.mlir:22060:28
  wire [31:0]     mult_inst214_result;	// matmul/matmul-hw.mlir:22030:28
  wire [31:0]     mult_inst213_result;	// matmul/matmul-hw.mlir:22000:28
  wire [31:0]     mult_inst212_result;	// matmul/matmul-hw.mlir:21970:28
  wire [31:0]     mult_inst211_result;	// matmul/matmul-hw.mlir:21940:28
  wire [31:0]     mult_inst210_result;	// matmul/matmul-hw.mlir:21910:28
  wire [31:0]     mult_inst209_result;	// matmul/matmul-hw.mlir:21880:28
  wire [31:0]     mult_inst208_result;	// matmul/matmul-hw.mlir:21850:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2216;	// matmul/matmul-hw.mlir:21845:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2217;	// matmul/matmul-hw.mlir:21844:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2218;	// matmul/matmul-hw.mlir:21843:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2219;	// matmul/matmul-hw.mlir:21842:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2220;	// matmul/matmul-hw.mlir:21841:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2221;	// matmul/matmul-hw.mlir:21840:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2222;	// matmul/matmul-hw.mlir:21839:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2223;	// matmul/matmul-hw.mlir:21838:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2224;	// matmul/matmul-hw.mlir:21837:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2225;	// matmul/matmul-hw.mlir:21836:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2226;	// matmul/matmul-hw.mlir:21835:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2227;	// matmul/matmul-hw.mlir:21834:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2228;	// matmul/matmul-hw.mlir:21833:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2229;	// matmul/matmul-hw.mlir:21832:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2230;	// matmul/matmul-hw.mlir:21831:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2231;	// matmul/matmul-hw.mlir:21830:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2232;	// matmul/matmul-hw.mlir:21829:36
  wire [31:0]     mult_inst207_result;	// matmul/matmul-hw.mlir:21690:28
  wire [31:0]     mult_inst206_result;	// matmul/matmul-hw.mlir:21660:28
  wire [31:0]     mult_inst205_result;	// matmul/matmul-hw.mlir:21630:28
  wire [31:0]     mult_inst204_result;	// matmul/matmul-hw.mlir:21600:28
  wire [31:0]     mult_inst203_result;	// matmul/matmul-hw.mlir:21570:28
  wire [31:0]     mult_inst202_result;	// matmul/matmul-hw.mlir:21540:28
  wire [31:0]     mult_inst201_result;	// matmul/matmul-hw.mlir:21510:28
  wire [31:0]     mult_inst200_result;	// matmul/matmul-hw.mlir:21480:28
  wire [31:0]     mult_inst199_result;	// matmul/matmul-hw.mlir:21450:28
  wire [31:0]     mult_inst198_result;	// matmul/matmul-hw.mlir:21420:28
  wire [31:0]     mult_inst197_result;	// matmul/matmul-hw.mlir:21390:28
  wire [31:0]     mult_inst196_result;	// matmul/matmul-hw.mlir:21360:28
  wire [31:0]     mult_inst195_result;	// matmul/matmul-hw.mlir:21330:28
  wire [31:0]     mult_inst194_result;	// matmul/matmul-hw.mlir:21300:28
  wire [31:0]     mult_inst193_result;	// matmul/matmul-hw.mlir:21270:28
  wire [31:0]     mult_inst192_result;	// matmul/matmul-hw.mlir:21240:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2233;	// matmul/matmul-hw.mlir:21235:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2234;	// matmul/matmul-hw.mlir:21234:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2235;	// matmul/matmul-hw.mlir:21233:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2236;	// matmul/matmul-hw.mlir:21232:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2237;	// matmul/matmul-hw.mlir:21231:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2238;	// matmul/matmul-hw.mlir:21230:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2239;	// matmul/matmul-hw.mlir:21229:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2240;	// matmul/matmul-hw.mlir:21228:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2241;	// matmul/matmul-hw.mlir:21227:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2242;	// matmul/matmul-hw.mlir:21226:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2243;	// matmul/matmul-hw.mlir:21225:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2244;	// matmul/matmul-hw.mlir:21224:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2245;	// matmul/matmul-hw.mlir:21223:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2246;	// matmul/matmul-hw.mlir:21222:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2247;	// matmul/matmul-hw.mlir:21221:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2248;	// matmul/matmul-hw.mlir:21220:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2249;	// matmul/matmul-hw.mlir:21219:36
  wire [31:0]     mult_inst191_result;	// matmul/matmul-hw.mlir:21095:28
  wire [31:0]     mult_inst190_result;	// matmul/matmul-hw.mlir:21065:28
  wire [31:0]     mult_inst189_result;	// matmul/matmul-hw.mlir:21035:28
  wire [31:0]     mult_inst188_result;	// matmul/matmul-hw.mlir:21005:28
  wire [31:0]     mult_inst187_result;	// matmul/matmul-hw.mlir:20975:28
  wire [31:0]     mult_inst186_result;	// matmul/matmul-hw.mlir:20945:28
  wire [31:0]     mult_inst185_result;	// matmul/matmul-hw.mlir:20915:28
  wire [31:0]     mult_inst184_result;	// matmul/matmul-hw.mlir:20885:28
  wire [31:0]     mult_inst183_result;	// matmul/matmul-hw.mlir:20855:28
  wire [31:0]     mult_inst182_result;	// matmul/matmul-hw.mlir:20825:28
  wire [31:0]     mult_inst181_result;	// matmul/matmul-hw.mlir:20795:28
  wire [31:0]     mult_inst180_result;	// matmul/matmul-hw.mlir:20765:28
  wire [31:0]     mult_inst179_result;	// matmul/matmul-hw.mlir:20735:28
  wire [31:0]     mult_inst178_result;	// matmul/matmul-hw.mlir:20705:28
  wire [31:0]     mult_inst177_result;	// matmul/matmul-hw.mlir:20675:28
  wire [31:0]     mult_inst176_result;	// matmul/matmul-hw.mlir:20645:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2250;	// matmul/matmul-hw.mlir:20640:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2251;	// matmul/matmul-hw.mlir:20639:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2252;	// matmul/matmul-hw.mlir:20638:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2253;	// matmul/matmul-hw.mlir:20637:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2254;	// matmul/matmul-hw.mlir:20636:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2255;	// matmul/matmul-hw.mlir:20635:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2256;	// matmul/matmul-hw.mlir:20634:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2257;	// matmul/matmul-hw.mlir:20633:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2258;	// matmul/matmul-hw.mlir:20632:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2259;	// matmul/matmul-hw.mlir:20631:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2260;	// matmul/matmul-hw.mlir:20630:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2261;	// matmul/matmul-hw.mlir:20629:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2262;	// matmul/matmul-hw.mlir:20628:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2263;	// matmul/matmul-hw.mlir:20627:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2264;	// matmul/matmul-hw.mlir:20626:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2265;	// matmul/matmul-hw.mlir:20625:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2266;	// matmul/matmul-hw.mlir:20624:36
  wire [31:0]     mult_inst175_result;	// matmul/matmul-hw.mlir:20500:28
  wire [31:0]     mult_inst174_result;	// matmul/matmul-hw.mlir:20470:28
  wire [31:0]     mult_inst173_result;	// matmul/matmul-hw.mlir:20440:28
  wire [31:0]     mult_inst172_result;	// matmul/matmul-hw.mlir:20410:28
  wire [31:0]     mult_inst171_result;	// matmul/matmul-hw.mlir:20380:28
  wire [31:0]     mult_inst170_result;	// matmul/matmul-hw.mlir:20350:28
  wire [31:0]     mult_inst169_result;	// matmul/matmul-hw.mlir:20320:28
  wire [31:0]     mult_inst168_result;	// matmul/matmul-hw.mlir:20290:28
  wire [31:0]     mult_inst167_result;	// matmul/matmul-hw.mlir:20260:28
  wire [31:0]     mult_inst166_result;	// matmul/matmul-hw.mlir:20230:28
  wire [31:0]     mult_inst165_result;	// matmul/matmul-hw.mlir:20200:28
  wire [31:0]     mult_inst164_result;	// matmul/matmul-hw.mlir:20170:28
  wire [31:0]     mult_inst163_result;	// matmul/matmul-hw.mlir:20140:28
  wire [31:0]     mult_inst162_result;	// matmul/matmul-hw.mlir:20110:28
  wire [31:0]     mult_inst161_result;	// matmul/matmul-hw.mlir:20080:28
  wire [31:0]     mult_inst160_result;	// matmul/matmul-hw.mlir:20050:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2267;	// matmul/matmul-hw.mlir:20045:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2268;	// matmul/matmul-hw.mlir:20044:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2269;	// matmul/matmul-hw.mlir:20043:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2270;	// matmul/matmul-hw.mlir:20042:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2271;	// matmul/matmul-hw.mlir:20041:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2272;	// matmul/matmul-hw.mlir:20040:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2273;	// matmul/matmul-hw.mlir:20039:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2274;	// matmul/matmul-hw.mlir:20038:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2275;	// matmul/matmul-hw.mlir:20037:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2276;	// matmul/matmul-hw.mlir:20036:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2277;	// matmul/matmul-hw.mlir:20035:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2278;	// matmul/matmul-hw.mlir:20034:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2279;	// matmul/matmul-hw.mlir:20033:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2280;	// matmul/matmul-hw.mlir:20032:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2281;	// matmul/matmul-hw.mlir:20031:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2282;	// matmul/matmul-hw.mlir:20030:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2283;	// matmul/matmul-hw.mlir:20029:36
  wire [31:0]     mult_inst159_result;	// matmul/matmul-hw.mlir:19905:28
  wire [31:0]     mult_inst158_result;	// matmul/matmul-hw.mlir:19875:28
  wire [31:0]     mult_inst157_result;	// matmul/matmul-hw.mlir:19845:28
  wire [31:0]     mult_inst156_result;	// matmul/matmul-hw.mlir:19815:28
  wire [31:0]     mult_inst155_result;	// matmul/matmul-hw.mlir:19785:28
  wire [31:0]     mult_inst154_result;	// matmul/matmul-hw.mlir:19755:28
  wire [31:0]     mult_inst153_result;	// matmul/matmul-hw.mlir:19725:28
  wire [31:0]     mult_inst152_result;	// matmul/matmul-hw.mlir:19695:28
  wire [31:0]     mult_inst151_result;	// matmul/matmul-hw.mlir:19665:28
  wire [31:0]     mult_inst150_result;	// matmul/matmul-hw.mlir:19635:28
  wire [31:0]     mult_inst149_result;	// matmul/matmul-hw.mlir:19605:28
  wire [31:0]     mult_inst148_result;	// matmul/matmul-hw.mlir:19575:28
  wire [31:0]     mult_inst147_result;	// matmul/matmul-hw.mlir:19545:28
  wire [31:0]     mult_inst146_result;	// matmul/matmul-hw.mlir:19515:28
  wire [31:0]     mult_inst145_result;	// matmul/matmul-hw.mlir:19485:28
  wire [31:0]     mult_inst144_result;	// matmul/matmul-hw.mlir:19455:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2284;	// matmul/matmul-hw.mlir:19450:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2285;	// matmul/matmul-hw.mlir:19449:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2286;	// matmul/matmul-hw.mlir:19448:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2287;	// matmul/matmul-hw.mlir:19447:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2288;	// matmul/matmul-hw.mlir:19446:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2289;	// matmul/matmul-hw.mlir:19445:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2290;	// matmul/matmul-hw.mlir:19444:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2291;	// matmul/matmul-hw.mlir:19443:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2292;	// matmul/matmul-hw.mlir:19442:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2293;	// matmul/matmul-hw.mlir:19441:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2294;	// matmul/matmul-hw.mlir:19440:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2295;	// matmul/matmul-hw.mlir:19439:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2296;	// matmul/matmul-hw.mlir:19438:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2297;	// matmul/matmul-hw.mlir:19437:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2298;	// matmul/matmul-hw.mlir:19436:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2299;	// matmul/matmul-hw.mlir:19435:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2300;	// matmul/matmul-hw.mlir:19434:36
  wire [31:0]     mult_inst143_result;	// matmul/matmul-hw.mlir:19310:28
  wire [31:0]     mult_inst142_result;	// matmul/matmul-hw.mlir:19280:28
  wire [31:0]     mult_inst141_result;	// matmul/matmul-hw.mlir:19250:28
  wire [31:0]     mult_inst140_result;	// matmul/matmul-hw.mlir:19220:28
  wire [31:0]     mult_inst139_result;	// matmul/matmul-hw.mlir:19190:28
  wire [31:0]     mult_inst138_result;	// matmul/matmul-hw.mlir:19160:28
  wire [31:0]     mult_inst137_result;	// matmul/matmul-hw.mlir:19130:28
  wire [31:0]     mult_inst136_result;	// matmul/matmul-hw.mlir:19100:28
  wire [31:0]     mult_inst135_result;	// matmul/matmul-hw.mlir:19070:28
  wire [31:0]     mult_inst134_result;	// matmul/matmul-hw.mlir:19040:28
  wire [31:0]     mult_inst133_result;	// matmul/matmul-hw.mlir:19010:28
  wire [31:0]     mult_inst132_result;	// matmul/matmul-hw.mlir:18980:28
  wire [31:0]     mult_inst131_result;	// matmul/matmul-hw.mlir:18950:28
  wire [31:0]     mult_inst130_result;	// matmul/matmul-hw.mlir:18920:28
  wire [31:0]     mult_inst129_result;	// matmul/matmul-hw.mlir:18890:28
  wire [31:0]     mult_inst128_result;	// matmul/matmul-hw.mlir:18860:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2301;	// matmul/matmul-hw.mlir:18855:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2302;	// matmul/matmul-hw.mlir:18854:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2303;	// matmul/matmul-hw.mlir:18853:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2304;	// matmul/matmul-hw.mlir:18852:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2305;	// matmul/matmul-hw.mlir:18851:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2306;	// matmul/matmul-hw.mlir:18850:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2307;	// matmul/matmul-hw.mlir:18849:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2308;	// matmul/matmul-hw.mlir:18848:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2309;	// matmul/matmul-hw.mlir:18847:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2310;	// matmul/matmul-hw.mlir:18846:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2311;	// matmul/matmul-hw.mlir:18845:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2312;	// matmul/matmul-hw.mlir:18844:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2313;	// matmul/matmul-hw.mlir:18843:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2314;	// matmul/matmul-hw.mlir:18842:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2315;	// matmul/matmul-hw.mlir:18841:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2316;	// matmul/matmul-hw.mlir:18840:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2317;	// matmul/matmul-hw.mlir:18839:36
  wire [31:0]     mult_inst127_result;	// matmul/matmul-hw.mlir:18715:28
  wire [31:0]     mult_inst126_result;	// matmul/matmul-hw.mlir:18685:28
  wire [31:0]     mult_inst125_result;	// matmul/matmul-hw.mlir:18655:28
  wire [31:0]     mult_inst124_result;	// matmul/matmul-hw.mlir:18625:28
  wire [31:0]     mult_inst123_result;	// matmul/matmul-hw.mlir:18595:28
  wire [31:0]     mult_inst122_result;	// matmul/matmul-hw.mlir:18565:28
  wire [31:0]     mult_inst121_result;	// matmul/matmul-hw.mlir:18535:28
  wire [31:0]     mult_inst120_result;	// matmul/matmul-hw.mlir:18505:28
  wire [31:0]     mult_inst119_result;	// matmul/matmul-hw.mlir:18475:28
  wire [31:0]     mult_inst118_result;	// matmul/matmul-hw.mlir:18445:28
  wire [31:0]     mult_inst117_result;	// matmul/matmul-hw.mlir:18415:28
  wire [31:0]     mult_inst116_result;	// matmul/matmul-hw.mlir:18385:28
  wire [31:0]     mult_inst115_result;	// matmul/matmul-hw.mlir:18355:28
  wire [31:0]     mult_inst114_result;	// matmul/matmul-hw.mlir:18325:28
  wire [31:0]     mult_inst113_result;	// matmul/matmul-hw.mlir:18295:28
  wire [31:0]     mult_inst112_result;	// matmul/matmul-hw.mlir:18265:28
  wire [31:0]     C_reg_bank16_p0_rd_data_2318;	// matmul/matmul-hw.mlir:18260:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2319;	// matmul/matmul-hw.mlir:18259:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2320;	// matmul/matmul-hw.mlir:18258:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2321;	// matmul/matmul-hw.mlir:18257:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2322;	// matmul/matmul-hw.mlir:18256:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2323;	// matmul/matmul-hw.mlir:18255:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2324;	// matmul/matmul-hw.mlir:18254:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2325;	// matmul/matmul-hw.mlir:18253:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2326;	// matmul/matmul-hw.mlir:18252:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2327;	// matmul/matmul-hw.mlir:18251:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2328;	// matmul/matmul-hw.mlir:18250:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2329;	// matmul/matmul-hw.mlir:18249:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2330;	// matmul/matmul-hw.mlir:18248:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2331;	// matmul/matmul-hw.mlir:18247:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2332;	// matmul/matmul-hw.mlir:18246:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2333;	// matmul/matmul-hw.mlir:18245:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2334;	// matmul/matmul-hw.mlir:18244:36
  wire [31:0]     mult_inst111_result;	// matmul/matmul-hw.mlir:18120:28
  wire [31:0]     mult_inst110_result;	// matmul/matmul-hw.mlir:18090:28
  wire [31:0]     mult_inst109_result;	// matmul/matmul-hw.mlir:18060:28
  wire [31:0]     mult_inst108_result;	// matmul/matmul-hw.mlir:18030:28
  wire [31:0]     mult_inst107_result;	// matmul/matmul-hw.mlir:18000:28
  wire [31:0]     mult_inst106_result;	// matmul/matmul-hw.mlir:17970:28
  wire [31:0]     mult_inst105_result;	// matmul/matmul-hw.mlir:17940:28
  wire [31:0]     mult_inst104_result;	// matmul/matmul-hw.mlir:17910:28
  wire [31:0]     mult_inst103_result;	// matmul/matmul-hw.mlir:17880:28
  wire [31:0]     mult_inst102_result;	// matmul/matmul-hw.mlir:17850:28
  wire [31:0]     mult_inst101_result;	// matmul/matmul-hw.mlir:17820:28
  wire [31:0]     mult_inst100_result;	// matmul/matmul-hw.mlir:17790:28
  wire [31:0]     mult_inst99_result;	// matmul/matmul-hw.mlir:17760:27
  wire [31:0]     mult_inst98_result;	// matmul/matmul-hw.mlir:17730:27
  wire [31:0]     mult_inst97_result;	// matmul/matmul-hw.mlir:17700:27
  wire [31:0]     mult_inst96_result;	// matmul/matmul-hw.mlir:17670:27
  wire [31:0]     C_reg_bank16_p0_rd_data_2335;	// matmul/matmul-hw.mlir:17665:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2336;	// matmul/matmul-hw.mlir:17664:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2337;	// matmul/matmul-hw.mlir:17663:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2338;	// matmul/matmul-hw.mlir:17662:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2339;	// matmul/matmul-hw.mlir:17661:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2340;	// matmul/matmul-hw.mlir:17660:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2341;	// matmul/matmul-hw.mlir:17659:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2342;	// matmul/matmul-hw.mlir:17658:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2343;	// matmul/matmul-hw.mlir:17657:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2344;	// matmul/matmul-hw.mlir:17656:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2345;	// matmul/matmul-hw.mlir:17655:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2346;	// matmul/matmul-hw.mlir:17654:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2347;	// matmul/matmul-hw.mlir:17653:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2348;	// matmul/matmul-hw.mlir:17652:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2349;	// matmul/matmul-hw.mlir:17651:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2350;	// matmul/matmul-hw.mlir:17650:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2351;	// matmul/matmul-hw.mlir:17649:36
  wire [31:0]     mult_inst95_result;	// matmul/matmul-hw.mlir:17525:27
  wire [31:0]     mult_inst94_result;	// matmul/matmul-hw.mlir:17495:27
  wire [31:0]     mult_inst93_result;	// matmul/matmul-hw.mlir:17465:27
  wire [31:0]     mult_inst92_result;	// matmul/matmul-hw.mlir:17435:27
  wire [31:0]     mult_inst91_result;	// matmul/matmul-hw.mlir:17405:27
  wire [31:0]     mult_inst90_result;	// matmul/matmul-hw.mlir:17375:27
  wire [31:0]     mult_inst89_result;	// matmul/matmul-hw.mlir:17345:27
  wire [31:0]     mult_inst88_result;	// matmul/matmul-hw.mlir:17315:27
  wire [31:0]     mult_inst87_result;	// matmul/matmul-hw.mlir:17285:27
  wire [31:0]     mult_inst86_result;	// matmul/matmul-hw.mlir:17255:27
  wire [31:0]     mult_inst85_result;	// matmul/matmul-hw.mlir:17225:27
  wire [31:0]     mult_inst84_result;	// matmul/matmul-hw.mlir:17195:27
  wire [31:0]     mult_inst83_result;	// matmul/matmul-hw.mlir:17165:27
  wire [31:0]     mult_inst82_result;	// matmul/matmul-hw.mlir:17135:27
  wire [31:0]     mult_inst81_result;	// matmul/matmul-hw.mlir:17105:27
  wire [31:0]     mult_inst80_result;	// matmul/matmul-hw.mlir:17075:27
  wire [31:0]     C_reg_bank16_p0_rd_data_2352;	// matmul/matmul-hw.mlir:17070:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2353;	// matmul/matmul-hw.mlir:17069:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2354;	// matmul/matmul-hw.mlir:17068:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2355;	// matmul/matmul-hw.mlir:17067:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2356;	// matmul/matmul-hw.mlir:17066:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2357;	// matmul/matmul-hw.mlir:17065:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2358;	// matmul/matmul-hw.mlir:17064:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2359;	// matmul/matmul-hw.mlir:17063:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2360;	// matmul/matmul-hw.mlir:17062:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2361;	// matmul/matmul-hw.mlir:17061:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2362;	// matmul/matmul-hw.mlir:17060:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2363;	// matmul/matmul-hw.mlir:17059:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2364;	// matmul/matmul-hw.mlir:17058:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2365;	// matmul/matmul-hw.mlir:17057:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2366;	// matmul/matmul-hw.mlir:17056:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2367;	// matmul/matmul-hw.mlir:17055:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2368;	// matmul/matmul-hw.mlir:17054:36
  wire [31:0]     mult_inst79_result;	// matmul/matmul-hw.mlir:16930:27
  wire [31:0]     mult_inst78_result;	// matmul/matmul-hw.mlir:16900:27
  wire [31:0]     mult_inst77_result;	// matmul/matmul-hw.mlir:16870:27
  wire [31:0]     mult_inst76_result;	// matmul/matmul-hw.mlir:16840:27
  wire [31:0]     mult_inst75_result;	// matmul/matmul-hw.mlir:16810:27
  wire [31:0]     mult_inst74_result;	// matmul/matmul-hw.mlir:16780:27
  wire [31:0]     mult_inst73_result;	// matmul/matmul-hw.mlir:16750:27
  wire [31:0]     mult_inst72_result;	// matmul/matmul-hw.mlir:16720:27
  wire [31:0]     mult_inst71_result;	// matmul/matmul-hw.mlir:16690:27
  wire [31:0]     mult_inst70_result;	// matmul/matmul-hw.mlir:16660:27
  wire [31:0]     mult_inst69_result;	// matmul/matmul-hw.mlir:16630:27
  wire [31:0]     mult_inst68_result;	// matmul/matmul-hw.mlir:16600:27
  wire [31:0]     mult_inst67_result;	// matmul/matmul-hw.mlir:16570:27
  wire [31:0]     mult_inst66_result;	// matmul/matmul-hw.mlir:16540:27
  wire [31:0]     mult_inst65_result;	// matmul/matmul-hw.mlir:16510:27
  wire [31:0]     mult_inst64_result;	// matmul/matmul-hw.mlir:16480:27
  wire [31:0]     C_reg_bank16_p0_rd_data_2369;	// matmul/matmul-hw.mlir:16475:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2370;	// matmul/matmul-hw.mlir:16474:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2371;	// matmul/matmul-hw.mlir:16473:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2372;	// matmul/matmul-hw.mlir:16472:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2373;	// matmul/matmul-hw.mlir:16471:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2374;	// matmul/matmul-hw.mlir:16470:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2375;	// matmul/matmul-hw.mlir:16469:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2376;	// matmul/matmul-hw.mlir:16468:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2377;	// matmul/matmul-hw.mlir:16467:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2378;	// matmul/matmul-hw.mlir:16466:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2379;	// matmul/matmul-hw.mlir:16465:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2380;	// matmul/matmul-hw.mlir:16464:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2381;	// matmul/matmul-hw.mlir:16463:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2382;	// matmul/matmul-hw.mlir:16462:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2383;	// matmul/matmul-hw.mlir:16461:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2384;	// matmul/matmul-hw.mlir:16460:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2385;	// matmul/matmul-hw.mlir:16459:36
  wire [31:0]     mult_inst63_result;	// matmul/matmul-hw.mlir:16335:27
  wire [31:0]     mult_inst62_result;	// matmul/matmul-hw.mlir:16305:27
  wire [31:0]     mult_inst61_result;	// matmul/matmul-hw.mlir:16275:27
  wire [31:0]     mult_inst60_result;	// matmul/matmul-hw.mlir:16245:27
  wire [31:0]     mult_inst59_result;	// matmul/matmul-hw.mlir:16215:27
  wire [31:0]     mult_inst58_result;	// matmul/matmul-hw.mlir:16185:27
  wire [31:0]     mult_inst57_result;	// matmul/matmul-hw.mlir:16155:27
  wire [31:0]     mult_inst56_result;	// matmul/matmul-hw.mlir:16125:27
  wire [31:0]     mult_inst55_result;	// matmul/matmul-hw.mlir:16095:27
  wire [31:0]     mult_inst54_result;	// matmul/matmul-hw.mlir:16065:27
  wire [31:0]     mult_inst53_result;	// matmul/matmul-hw.mlir:16035:27
  wire [31:0]     mult_inst52_result;	// matmul/matmul-hw.mlir:16005:27
  wire [31:0]     mult_inst51_result;	// matmul/matmul-hw.mlir:15975:27
  wire [31:0]     mult_inst50_result;	// matmul/matmul-hw.mlir:15945:27
  wire [31:0]     mult_inst49_result;	// matmul/matmul-hw.mlir:15915:27
  wire [31:0]     mult_inst48_result;	// matmul/matmul-hw.mlir:15885:27
  wire [31:0]     C_reg_bank16_p0_rd_data_2386;	// matmul/matmul-hw.mlir:15880:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2387;	// matmul/matmul-hw.mlir:15879:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2388;	// matmul/matmul-hw.mlir:15878:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2389;	// matmul/matmul-hw.mlir:15877:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2390;	// matmul/matmul-hw.mlir:15876:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2391;	// matmul/matmul-hw.mlir:15875:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2392;	// matmul/matmul-hw.mlir:15874:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2393;	// matmul/matmul-hw.mlir:15873:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2394;	// matmul/matmul-hw.mlir:15872:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2395;	// matmul/matmul-hw.mlir:15871:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2396;	// matmul/matmul-hw.mlir:15870:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2397;	// matmul/matmul-hw.mlir:15869:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2398;	// matmul/matmul-hw.mlir:15868:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2399;	// matmul/matmul-hw.mlir:15867:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2400;	// matmul/matmul-hw.mlir:15866:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2401;	// matmul/matmul-hw.mlir:15865:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2402;	// matmul/matmul-hw.mlir:15864:36
  wire [31:0]     mult_inst47_result;	// matmul/matmul-hw.mlir:15740:27
  wire [31:0]     mult_inst46_result;	// matmul/matmul-hw.mlir:15710:27
  wire [31:0]     mult_inst45_result;	// matmul/matmul-hw.mlir:15680:27
  wire [31:0]     mult_inst44_result;	// matmul/matmul-hw.mlir:15650:27
  wire [31:0]     mult_inst43_result;	// matmul/matmul-hw.mlir:15620:27
  wire [31:0]     mult_inst42_result;	// matmul/matmul-hw.mlir:15590:27
  wire [31:0]     mult_inst41_result;	// matmul/matmul-hw.mlir:15560:27
  wire [31:0]     mult_inst40_result;	// matmul/matmul-hw.mlir:15530:27
  wire [31:0]     mult_inst39_result;	// matmul/matmul-hw.mlir:15500:27
  wire [31:0]     mult_inst38_result;	// matmul/matmul-hw.mlir:15470:27
  wire [31:0]     mult_inst37_result;	// matmul/matmul-hw.mlir:15440:27
  wire [31:0]     mult_inst36_result;	// matmul/matmul-hw.mlir:15410:27
  wire [31:0]     mult_inst35_result;	// matmul/matmul-hw.mlir:15380:27
  wire [31:0]     mult_inst34_result;	// matmul/matmul-hw.mlir:15350:27
  wire [31:0]     mult_inst33_result;	// matmul/matmul-hw.mlir:15320:27
  wire [31:0]     mult_inst32_result;	// matmul/matmul-hw.mlir:15290:27
  wire [31:0]     C_reg_bank16_p0_rd_data_2403;	// matmul/matmul-hw.mlir:15285:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2404;	// matmul/matmul-hw.mlir:15284:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2405;	// matmul/matmul-hw.mlir:15283:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2406;	// matmul/matmul-hw.mlir:15282:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2407;	// matmul/matmul-hw.mlir:15281:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2408;	// matmul/matmul-hw.mlir:15280:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2409;	// matmul/matmul-hw.mlir:15279:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2410;	// matmul/matmul-hw.mlir:15278:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2411;	// matmul/matmul-hw.mlir:15277:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2412;	// matmul/matmul-hw.mlir:15276:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2413;	// matmul/matmul-hw.mlir:15275:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2414;	// matmul/matmul-hw.mlir:15274:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2415;	// matmul/matmul-hw.mlir:15273:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2416;	// matmul/matmul-hw.mlir:15272:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2417;	// matmul/matmul-hw.mlir:15271:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2418;	// matmul/matmul-hw.mlir:15270:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2419;	// matmul/matmul-hw.mlir:15269:36
  wire [31:0]     mult_inst31_result;	// matmul/matmul-hw.mlir:15145:27
  wire [31:0]     mult_inst30_result;	// matmul/matmul-hw.mlir:15115:27
  wire [31:0]     mult_inst29_result;	// matmul/matmul-hw.mlir:15085:27
  wire [31:0]     mult_inst28_result;	// matmul/matmul-hw.mlir:15055:27
  wire [31:0]     mult_inst27_result;	// matmul/matmul-hw.mlir:15025:27
  wire [31:0]     mult_inst26_result;	// matmul/matmul-hw.mlir:14995:27
  wire [31:0]     mult_inst25_result;	// matmul/matmul-hw.mlir:14965:27
  wire [31:0]     mult_inst24_result;	// matmul/matmul-hw.mlir:14935:27
  wire [31:0]     mult_inst23_result;	// matmul/matmul-hw.mlir:14905:27
  wire [31:0]     mult_inst22_result;	// matmul/matmul-hw.mlir:14875:27
  wire [31:0]     mult_inst21_result;	// matmul/matmul-hw.mlir:14845:27
  wire [31:0]     mult_inst20_result;	// matmul/matmul-hw.mlir:14815:27
  wire [31:0]     mult_inst19_result;	// matmul/matmul-hw.mlir:14785:27
  wire [31:0]     mult_inst18_result;	// matmul/matmul-hw.mlir:14755:27
  wire [31:0]     mult_inst17_result;	// matmul/matmul-hw.mlir:14725:27
  wire [31:0]     mult_inst16_result;	// matmul/matmul-hw.mlir:14695:27
  wire [31:0]     C_reg_bank16_p0_rd_data_2420;	// matmul/matmul-hw.mlir:14690:37
  wire [31:0]     C_reg_bank15_p0_rd_data_2421;	// matmul/matmul-hw.mlir:14689:37
  wire [31:0]     C_reg_bank14_p0_rd_data_2422;	// matmul/matmul-hw.mlir:14688:37
  wire [31:0]     C_reg_bank13_p0_rd_data_2423;	// matmul/matmul-hw.mlir:14687:37
  wire [31:0]     C_reg_bank12_p0_rd_data_2424;	// matmul/matmul-hw.mlir:14686:37
  wire [31:0]     C_reg_bank11_p0_rd_data_2425;	// matmul/matmul-hw.mlir:14685:37
  wire [31:0]     C_reg_bank10_p0_rd_data_2426;	// matmul/matmul-hw.mlir:14684:37
  wire [31:0]     C_reg_bank9_p0_rd_data_2427;	// matmul/matmul-hw.mlir:14683:36
  wire [31:0]     C_reg_bank8_p0_rd_data_2428;	// matmul/matmul-hw.mlir:14682:36
  wire [31:0]     C_reg_bank7_p0_rd_data_2429;	// matmul/matmul-hw.mlir:14681:36
  wire [31:0]     C_reg_bank6_p0_rd_data_2430;	// matmul/matmul-hw.mlir:14680:36
  wire [31:0]     C_reg_bank5_p0_rd_data_2431;	// matmul/matmul-hw.mlir:14679:36
  wire [31:0]     C_reg_bank4_p0_rd_data_2432;	// matmul/matmul-hw.mlir:14678:36
  wire [31:0]     C_reg_bank3_p0_rd_data_2433;	// matmul/matmul-hw.mlir:14677:36
  wire [31:0]     C_reg_bank2_p0_rd_data_2434;	// matmul/matmul-hw.mlir:14676:36
  wire [31:0]     C_reg_bank1_p0_rd_data_2435;	// matmul/matmul-hw.mlir:14675:36
  wire [31:0]     C_reg_bank0_p0_rd_data_2436;	// matmul/matmul-hw.mlir:14674:36
  wire [31:0]     mult_inst15_result;	// matmul/matmul-hw.mlir:14558:27
  wire [31:0]     mult_inst14_result;	// matmul/matmul-hw.mlir:14536:27
  wire [31:0]     mult_inst13_result;	// matmul/matmul-hw.mlir:14514:27
  wire [31:0]     mult_inst12_result;	// matmul/matmul-hw.mlir:14492:27
  wire [31:0]     mult_inst11_result;	// matmul/matmul-hw.mlir:14470:27
  wire [31:0]     mult_inst10_result;	// matmul/matmul-hw.mlir:14448:27
  wire [31:0]     mult_inst9_result;	// matmul/matmul-hw.mlir:14426:26
  wire [31:0]     mult_inst8_result;	// matmul/matmul-hw.mlir:14404:26
  wire [31:0]     mult_inst7_result;	// matmul/matmul-hw.mlir:14382:26
  wire [31:0]     mult_inst6_result;	// matmul/matmul-hw.mlir:14360:26
  wire [31:0]     mult_inst5_result;	// matmul/matmul-hw.mlir:14338:26
  wire [31:0]     mult_inst4_result;	// matmul/matmul-hw.mlir:14316:26
  wire [31:0]     mult_inst3_result;	// matmul/matmul-hw.mlir:14294:26
  wire [31:0]     mult_inst2_result;	// matmul/matmul-hw.mlir:14272:26
  wire [31:0]     mult_inst1_result;	// matmul/matmul-hw.mlir:14250:26
  wire [31:0]     mult_inst0_result;	// matmul/matmul-hw.mlir:14228:26
  wire [31:0]     C_reg_bank16_p0_rd_data_2437;	// matmul/matmul-hw.mlir:14223:32
  wire [31:0]     C_reg_bank15_p0_rd_data_2438;	// matmul/matmul-hw.mlir:14222:32
  wire [31:0]     C_reg_bank14_p0_rd_data_2439;	// matmul/matmul-hw.mlir:14221:32
  wire [31:0]     C_reg_bank13_p0_rd_data_2440;	// matmul/matmul-hw.mlir:14220:32
  wire [31:0]     C_reg_bank12_p0_rd_data_2441;	// matmul/matmul-hw.mlir:14219:32
  wire [31:0]     C_reg_bank11_p0_rd_data_2442;	// matmul/matmul-hw.mlir:14218:32
  wire [31:0]     C_reg_bank10_p0_rd_data_2443;	// matmul/matmul-hw.mlir:14217:32
  wire [31:0]     C_reg_bank9_p0_rd_data_2444;	// matmul/matmul-hw.mlir:14216:31
  wire [31:0]     C_reg_bank8_p0_rd_data_2445;	// matmul/matmul-hw.mlir:14215:31
  wire [31:0]     C_reg_bank7_p0_rd_data_2446;	// matmul/matmul-hw.mlir:14214:31
  wire [31:0]     C_reg_bank6_p0_rd_data_2447;	// matmul/matmul-hw.mlir:14213:31
  wire [31:0]     C_reg_bank5_p0_rd_data_2448;	// matmul/matmul-hw.mlir:14212:31
  wire [31:0]     C_reg_bank4_p0_rd_data_2449;	// matmul/matmul-hw.mlir:14211:31
  wire [31:0]     C_reg_bank3_p0_rd_data_2450;	// matmul/matmul-hw.mlir:14210:31
  wire [31:0]     C_reg_bank2_p0_rd_data_2451;	// matmul/matmul-hw.mlir:14209:31
  wire [31:0]     C_reg_bank1_p0_rd_data_2452;	// matmul/matmul-hw.mlir:14208:31
  wire [31:0]     C_reg_bank0_p0_rd_data_2453;	// matmul/matmul-hw.mlir:14207:31
  wire [31:0]     A_reg_bank255_p0_rd_data;	// matmul/matmul-hw.mlir:12470:33
  wire [31:0]     A_reg_bank254_p0_rd_data;	// matmul/matmul-hw.mlir:12469:33
  wire [31:0]     A_reg_bank253_p0_rd_data;	// matmul/matmul-hw.mlir:12468:33
  wire [31:0]     A_reg_bank252_p0_rd_data;	// matmul/matmul-hw.mlir:12467:33
  wire [31:0]     A_reg_bank251_p0_rd_data;	// matmul/matmul-hw.mlir:12466:33
  wire [31:0]     A_reg_bank250_p0_rd_data;	// matmul/matmul-hw.mlir:12465:33
  wire [31:0]     A_reg_bank249_p0_rd_data;	// matmul/matmul-hw.mlir:12464:33
  wire [31:0]     A_reg_bank248_p0_rd_data;	// matmul/matmul-hw.mlir:12463:33
  wire [31:0]     A_reg_bank247_p0_rd_data;	// matmul/matmul-hw.mlir:12462:33
  wire [31:0]     A_reg_bank246_p0_rd_data;	// matmul/matmul-hw.mlir:12461:33
  wire [31:0]     A_reg_bank245_p0_rd_data;	// matmul/matmul-hw.mlir:12460:33
  wire [31:0]     A_reg_bank244_p0_rd_data;	// matmul/matmul-hw.mlir:12459:33
  wire [31:0]     A_reg_bank243_p0_rd_data;	// matmul/matmul-hw.mlir:12458:33
  wire [31:0]     A_reg_bank242_p0_rd_data;	// matmul/matmul-hw.mlir:12457:33
  wire [31:0]     A_reg_bank241_p0_rd_data;	// matmul/matmul-hw.mlir:12456:33
  wire [31:0]     A_reg_bank240_p0_rd_data;	// matmul/matmul-hw.mlir:12455:33
  wire [31:0]     A_reg_bank239_p0_rd_data;	// matmul/matmul-hw.mlir:12454:33
  wire [31:0]     A_reg_bank238_p0_rd_data;	// matmul/matmul-hw.mlir:12453:33
  wire [31:0]     A_reg_bank237_p0_rd_data;	// matmul/matmul-hw.mlir:12452:33
  wire [31:0]     A_reg_bank236_p0_rd_data;	// matmul/matmul-hw.mlir:12451:33
  wire [31:0]     A_reg_bank235_p0_rd_data;	// matmul/matmul-hw.mlir:12450:33
  wire [31:0]     A_reg_bank234_p0_rd_data;	// matmul/matmul-hw.mlir:12449:33
  wire [31:0]     A_reg_bank233_p0_rd_data;	// matmul/matmul-hw.mlir:12448:33
  wire [31:0]     A_reg_bank232_p0_rd_data;	// matmul/matmul-hw.mlir:12447:33
  wire [31:0]     A_reg_bank231_p0_rd_data;	// matmul/matmul-hw.mlir:12446:33
  wire [31:0]     A_reg_bank230_p0_rd_data;	// matmul/matmul-hw.mlir:12445:33
  wire [31:0]     A_reg_bank229_p0_rd_data;	// matmul/matmul-hw.mlir:12444:33
  wire [31:0]     A_reg_bank228_p0_rd_data;	// matmul/matmul-hw.mlir:12443:33
  wire [31:0]     A_reg_bank227_p0_rd_data;	// matmul/matmul-hw.mlir:12442:33
  wire [31:0]     A_reg_bank226_p0_rd_data;	// matmul/matmul-hw.mlir:12441:33
  wire [31:0]     A_reg_bank225_p0_rd_data;	// matmul/matmul-hw.mlir:12440:33
  wire [31:0]     A_reg_bank224_p0_rd_data;	// matmul/matmul-hw.mlir:12439:33
  wire [31:0]     A_reg_bank223_p0_rd_data;	// matmul/matmul-hw.mlir:12438:33
  wire [31:0]     A_reg_bank222_p0_rd_data;	// matmul/matmul-hw.mlir:12437:33
  wire [31:0]     A_reg_bank221_p0_rd_data;	// matmul/matmul-hw.mlir:12436:33
  wire [31:0]     A_reg_bank220_p0_rd_data;	// matmul/matmul-hw.mlir:12435:33
  wire [31:0]     A_reg_bank219_p0_rd_data;	// matmul/matmul-hw.mlir:12434:33
  wire [31:0]     A_reg_bank218_p0_rd_data;	// matmul/matmul-hw.mlir:12433:33
  wire [31:0]     A_reg_bank217_p0_rd_data;	// matmul/matmul-hw.mlir:12432:33
  wire [31:0]     A_reg_bank216_p0_rd_data;	// matmul/matmul-hw.mlir:12431:33
  wire [31:0]     A_reg_bank215_p0_rd_data;	// matmul/matmul-hw.mlir:12430:33
  wire [31:0]     A_reg_bank214_p0_rd_data;	// matmul/matmul-hw.mlir:12429:33
  wire [31:0]     A_reg_bank213_p0_rd_data;	// matmul/matmul-hw.mlir:12428:33
  wire [31:0]     A_reg_bank212_p0_rd_data;	// matmul/matmul-hw.mlir:12427:33
  wire [31:0]     A_reg_bank211_p0_rd_data;	// matmul/matmul-hw.mlir:12426:33
  wire [31:0]     A_reg_bank210_p0_rd_data;	// matmul/matmul-hw.mlir:12425:33
  wire [31:0]     A_reg_bank209_p0_rd_data;	// matmul/matmul-hw.mlir:12424:33
  wire [31:0]     A_reg_bank208_p0_rd_data;	// matmul/matmul-hw.mlir:12423:33
  wire [31:0]     A_reg_bank207_p0_rd_data;	// matmul/matmul-hw.mlir:12422:33
  wire [31:0]     A_reg_bank206_p0_rd_data;	// matmul/matmul-hw.mlir:12421:33
  wire [31:0]     A_reg_bank205_p0_rd_data;	// matmul/matmul-hw.mlir:12420:33
  wire [31:0]     A_reg_bank204_p0_rd_data;	// matmul/matmul-hw.mlir:12419:33
  wire [31:0]     A_reg_bank203_p0_rd_data;	// matmul/matmul-hw.mlir:12418:33
  wire [31:0]     A_reg_bank202_p0_rd_data;	// matmul/matmul-hw.mlir:12417:33
  wire [31:0]     A_reg_bank201_p0_rd_data;	// matmul/matmul-hw.mlir:12416:33
  wire [31:0]     A_reg_bank200_p0_rd_data;	// matmul/matmul-hw.mlir:12415:33
  wire [31:0]     A_reg_bank199_p0_rd_data;	// matmul/matmul-hw.mlir:12414:33
  wire [31:0]     A_reg_bank198_p0_rd_data;	// matmul/matmul-hw.mlir:12413:33
  wire [31:0]     A_reg_bank197_p0_rd_data;	// matmul/matmul-hw.mlir:12412:33
  wire [31:0]     A_reg_bank196_p0_rd_data;	// matmul/matmul-hw.mlir:12411:33
  wire [31:0]     A_reg_bank195_p0_rd_data;	// matmul/matmul-hw.mlir:12410:33
  wire [31:0]     A_reg_bank194_p0_rd_data;	// matmul/matmul-hw.mlir:12409:33
  wire [31:0]     A_reg_bank193_p0_rd_data;	// matmul/matmul-hw.mlir:12408:33
  wire [31:0]     A_reg_bank192_p0_rd_data;	// matmul/matmul-hw.mlir:12407:33
  wire [31:0]     A_reg_bank191_p0_rd_data;	// matmul/matmul-hw.mlir:12406:33
  wire [31:0]     A_reg_bank190_p0_rd_data;	// matmul/matmul-hw.mlir:12405:33
  wire [31:0]     A_reg_bank189_p0_rd_data;	// matmul/matmul-hw.mlir:12404:33
  wire [31:0]     A_reg_bank188_p0_rd_data;	// matmul/matmul-hw.mlir:12403:33
  wire [31:0]     A_reg_bank187_p0_rd_data;	// matmul/matmul-hw.mlir:12402:33
  wire [31:0]     A_reg_bank186_p0_rd_data;	// matmul/matmul-hw.mlir:12401:33
  wire [31:0]     A_reg_bank185_p0_rd_data;	// matmul/matmul-hw.mlir:12400:33
  wire [31:0]     A_reg_bank184_p0_rd_data;	// matmul/matmul-hw.mlir:12399:33
  wire [31:0]     A_reg_bank183_p0_rd_data;	// matmul/matmul-hw.mlir:12398:33
  wire [31:0]     A_reg_bank182_p0_rd_data;	// matmul/matmul-hw.mlir:12397:33
  wire [31:0]     A_reg_bank181_p0_rd_data;	// matmul/matmul-hw.mlir:12396:33
  wire [31:0]     A_reg_bank180_p0_rd_data;	// matmul/matmul-hw.mlir:12395:33
  wire [31:0]     A_reg_bank179_p0_rd_data;	// matmul/matmul-hw.mlir:12394:33
  wire [31:0]     A_reg_bank178_p0_rd_data;	// matmul/matmul-hw.mlir:12393:33
  wire [31:0]     A_reg_bank177_p0_rd_data;	// matmul/matmul-hw.mlir:12392:33
  wire [31:0]     A_reg_bank176_p0_rd_data;	// matmul/matmul-hw.mlir:12391:33
  wire [31:0]     A_reg_bank175_p0_rd_data;	// matmul/matmul-hw.mlir:12390:33
  wire [31:0]     A_reg_bank174_p0_rd_data;	// matmul/matmul-hw.mlir:12389:33
  wire [31:0]     A_reg_bank173_p0_rd_data;	// matmul/matmul-hw.mlir:12388:33
  wire [31:0]     A_reg_bank172_p0_rd_data;	// matmul/matmul-hw.mlir:12387:33
  wire [31:0]     A_reg_bank171_p0_rd_data;	// matmul/matmul-hw.mlir:12386:33
  wire [31:0]     A_reg_bank170_p0_rd_data;	// matmul/matmul-hw.mlir:12385:33
  wire [31:0]     A_reg_bank169_p0_rd_data;	// matmul/matmul-hw.mlir:12384:33
  wire [31:0]     A_reg_bank168_p0_rd_data;	// matmul/matmul-hw.mlir:12383:33
  wire [31:0]     A_reg_bank167_p0_rd_data;	// matmul/matmul-hw.mlir:12382:33
  wire [31:0]     A_reg_bank166_p0_rd_data;	// matmul/matmul-hw.mlir:12381:33
  wire [31:0]     A_reg_bank165_p0_rd_data;	// matmul/matmul-hw.mlir:12380:33
  wire [31:0]     A_reg_bank164_p0_rd_data;	// matmul/matmul-hw.mlir:12379:33
  wire [31:0]     A_reg_bank163_p0_rd_data;	// matmul/matmul-hw.mlir:12378:33
  wire [31:0]     A_reg_bank162_p0_rd_data;	// matmul/matmul-hw.mlir:12377:33
  wire [31:0]     A_reg_bank161_p0_rd_data;	// matmul/matmul-hw.mlir:12376:33
  wire [31:0]     A_reg_bank160_p0_rd_data;	// matmul/matmul-hw.mlir:12375:33
  wire [31:0]     A_reg_bank159_p0_rd_data;	// matmul/matmul-hw.mlir:12374:33
  wire [31:0]     A_reg_bank158_p0_rd_data;	// matmul/matmul-hw.mlir:12373:33
  wire [31:0]     A_reg_bank157_p0_rd_data;	// matmul/matmul-hw.mlir:12372:33
  wire [31:0]     A_reg_bank156_p0_rd_data;	// matmul/matmul-hw.mlir:12371:33
  wire [31:0]     A_reg_bank155_p0_rd_data;	// matmul/matmul-hw.mlir:12370:33
  wire [31:0]     A_reg_bank154_p0_rd_data;	// matmul/matmul-hw.mlir:12369:33
  wire [31:0]     A_reg_bank153_p0_rd_data;	// matmul/matmul-hw.mlir:12368:33
  wire [31:0]     A_reg_bank152_p0_rd_data;	// matmul/matmul-hw.mlir:12367:33
  wire [31:0]     A_reg_bank151_p0_rd_data;	// matmul/matmul-hw.mlir:12366:33
  wire [31:0]     A_reg_bank150_p0_rd_data;	// matmul/matmul-hw.mlir:12365:33
  wire [31:0]     A_reg_bank149_p0_rd_data;	// matmul/matmul-hw.mlir:12364:33
  wire [31:0]     A_reg_bank148_p0_rd_data;	// matmul/matmul-hw.mlir:12363:33
  wire [31:0]     A_reg_bank147_p0_rd_data;	// matmul/matmul-hw.mlir:12362:33
  wire [31:0]     A_reg_bank146_p0_rd_data;	// matmul/matmul-hw.mlir:12361:33
  wire [31:0]     A_reg_bank145_p0_rd_data;	// matmul/matmul-hw.mlir:12360:33
  wire [31:0]     A_reg_bank144_p0_rd_data;	// matmul/matmul-hw.mlir:12359:33
  wire [31:0]     A_reg_bank143_p0_rd_data;	// matmul/matmul-hw.mlir:12358:33
  wire [31:0]     A_reg_bank142_p0_rd_data;	// matmul/matmul-hw.mlir:12357:33
  wire [31:0]     A_reg_bank141_p0_rd_data;	// matmul/matmul-hw.mlir:12356:33
  wire [31:0]     A_reg_bank140_p0_rd_data;	// matmul/matmul-hw.mlir:12355:33
  wire [31:0]     A_reg_bank139_p0_rd_data;	// matmul/matmul-hw.mlir:12354:33
  wire [31:0]     A_reg_bank138_p0_rd_data;	// matmul/matmul-hw.mlir:12353:33
  wire [31:0]     A_reg_bank137_p0_rd_data;	// matmul/matmul-hw.mlir:12352:33
  wire [31:0]     A_reg_bank136_p0_rd_data;	// matmul/matmul-hw.mlir:12351:33
  wire [31:0]     A_reg_bank135_p0_rd_data;	// matmul/matmul-hw.mlir:12350:33
  wire [31:0]     A_reg_bank134_p0_rd_data;	// matmul/matmul-hw.mlir:12349:33
  wire [31:0]     A_reg_bank133_p0_rd_data;	// matmul/matmul-hw.mlir:12348:33
  wire [31:0]     A_reg_bank132_p0_rd_data;	// matmul/matmul-hw.mlir:12347:33
  wire [31:0]     A_reg_bank131_p0_rd_data;	// matmul/matmul-hw.mlir:12346:33
  wire [31:0]     A_reg_bank130_p0_rd_data;	// matmul/matmul-hw.mlir:12345:33
  wire [31:0]     A_reg_bank129_p0_rd_data;	// matmul/matmul-hw.mlir:12344:33
  wire [31:0]     A_reg_bank128_p0_rd_data;	// matmul/matmul-hw.mlir:12343:33
  wire [31:0]     A_reg_bank127_p0_rd_data;	// matmul/matmul-hw.mlir:12342:33
  wire [31:0]     A_reg_bank126_p0_rd_data;	// matmul/matmul-hw.mlir:12341:33
  wire [31:0]     A_reg_bank125_p0_rd_data;	// matmul/matmul-hw.mlir:12340:33
  wire [31:0]     A_reg_bank124_p0_rd_data;	// matmul/matmul-hw.mlir:12339:33
  wire [31:0]     A_reg_bank123_p0_rd_data;	// matmul/matmul-hw.mlir:12338:33
  wire [31:0]     A_reg_bank122_p0_rd_data;	// matmul/matmul-hw.mlir:12337:33
  wire [31:0]     A_reg_bank121_p0_rd_data;	// matmul/matmul-hw.mlir:12336:33
  wire [31:0]     A_reg_bank120_p0_rd_data;	// matmul/matmul-hw.mlir:12335:33
  wire [31:0]     A_reg_bank119_p0_rd_data;	// matmul/matmul-hw.mlir:12334:33
  wire [31:0]     A_reg_bank118_p0_rd_data;	// matmul/matmul-hw.mlir:12333:33
  wire [31:0]     A_reg_bank117_p0_rd_data;	// matmul/matmul-hw.mlir:12332:33
  wire [31:0]     A_reg_bank116_p0_rd_data;	// matmul/matmul-hw.mlir:12331:33
  wire [31:0]     A_reg_bank115_p0_rd_data;	// matmul/matmul-hw.mlir:12330:33
  wire [31:0]     A_reg_bank114_p0_rd_data;	// matmul/matmul-hw.mlir:12329:33
  wire [31:0]     A_reg_bank113_p0_rd_data;	// matmul/matmul-hw.mlir:12328:33
  wire [31:0]     A_reg_bank112_p0_rd_data;	// matmul/matmul-hw.mlir:12327:33
  wire [31:0]     A_reg_bank111_p0_rd_data;	// matmul/matmul-hw.mlir:12326:33
  wire [31:0]     A_reg_bank110_p0_rd_data;	// matmul/matmul-hw.mlir:12325:33
  wire [31:0]     A_reg_bank109_p0_rd_data;	// matmul/matmul-hw.mlir:12324:33
  wire [31:0]     A_reg_bank108_p0_rd_data;	// matmul/matmul-hw.mlir:12323:33
  wire [31:0]     A_reg_bank107_p0_rd_data;	// matmul/matmul-hw.mlir:12322:33
  wire [31:0]     A_reg_bank106_p0_rd_data;	// matmul/matmul-hw.mlir:12321:33
  wire [31:0]     A_reg_bank105_p0_rd_data;	// matmul/matmul-hw.mlir:12320:33
  wire [31:0]     A_reg_bank104_p0_rd_data;	// matmul/matmul-hw.mlir:12319:33
  wire [31:0]     A_reg_bank103_p0_rd_data;	// matmul/matmul-hw.mlir:12318:33
  wire [31:0]     A_reg_bank102_p0_rd_data;	// matmul/matmul-hw.mlir:12317:33
  wire [31:0]     A_reg_bank101_p0_rd_data;	// matmul/matmul-hw.mlir:12316:33
  wire [31:0]     A_reg_bank100_p0_rd_data;	// matmul/matmul-hw.mlir:12315:33
  wire [31:0]     A_reg_bank99_p0_rd_data;	// matmul/matmul-hw.mlir:12314:32
  wire [31:0]     A_reg_bank98_p0_rd_data;	// matmul/matmul-hw.mlir:12313:32
  wire [31:0]     A_reg_bank97_p0_rd_data;	// matmul/matmul-hw.mlir:12312:32
  wire [31:0]     A_reg_bank96_p0_rd_data;	// matmul/matmul-hw.mlir:12311:32
  wire [31:0]     A_reg_bank95_p0_rd_data;	// matmul/matmul-hw.mlir:12310:32
  wire [31:0]     A_reg_bank94_p0_rd_data;	// matmul/matmul-hw.mlir:12309:32
  wire [31:0]     A_reg_bank93_p0_rd_data;	// matmul/matmul-hw.mlir:12308:32
  wire [31:0]     A_reg_bank92_p0_rd_data;	// matmul/matmul-hw.mlir:12307:32
  wire [31:0]     A_reg_bank91_p0_rd_data;	// matmul/matmul-hw.mlir:12306:32
  wire [31:0]     A_reg_bank90_p0_rd_data;	// matmul/matmul-hw.mlir:12305:32
  wire [31:0]     A_reg_bank89_p0_rd_data;	// matmul/matmul-hw.mlir:12304:32
  wire [31:0]     A_reg_bank88_p0_rd_data;	// matmul/matmul-hw.mlir:12303:32
  wire [31:0]     A_reg_bank87_p0_rd_data;	// matmul/matmul-hw.mlir:12302:32
  wire [31:0]     A_reg_bank86_p0_rd_data;	// matmul/matmul-hw.mlir:12301:32
  wire [31:0]     A_reg_bank85_p0_rd_data;	// matmul/matmul-hw.mlir:12300:32
  wire [31:0]     A_reg_bank84_p0_rd_data;	// matmul/matmul-hw.mlir:12299:32
  wire [31:0]     A_reg_bank83_p0_rd_data;	// matmul/matmul-hw.mlir:12298:32
  wire [31:0]     A_reg_bank82_p0_rd_data;	// matmul/matmul-hw.mlir:12297:32
  wire [31:0]     A_reg_bank81_p0_rd_data;	// matmul/matmul-hw.mlir:12296:32
  wire [31:0]     A_reg_bank80_p0_rd_data;	// matmul/matmul-hw.mlir:12295:32
  wire [31:0]     A_reg_bank79_p0_rd_data;	// matmul/matmul-hw.mlir:12294:32
  wire [31:0]     A_reg_bank78_p0_rd_data;	// matmul/matmul-hw.mlir:12293:32
  wire [31:0]     A_reg_bank77_p0_rd_data;	// matmul/matmul-hw.mlir:12292:32
  wire [31:0]     A_reg_bank76_p0_rd_data;	// matmul/matmul-hw.mlir:12291:32
  wire [31:0]     A_reg_bank75_p0_rd_data;	// matmul/matmul-hw.mlir:12290:32
  wire [31:0]     A_reg_bank74_p0_rd_data;	// matmul/matmul-hw.mlir:12289:32
  wire [31:0]     A_reg_bank73_p0_rd_data;	// matmul/matmul-hw.mlir:12288:32
  wire [31:0]     A_reg_bank72_p0_rd_data;	// matmul/matmul-hw.mlir:12287:32
  wire [31:0]     A_reg_bank71_p0_rd_data;	// matmul/matmul-hw.mlir:12286:32
  wire [31:0]     A_reg_bank70_p0_rd_data;	// matmul/matmul-hw.mlir:12285:32
  wire [31:0]     A_reg_bank69_p0_rd_data;	// matmul/matmul-hw.mlir:12284:32
  wire [31:0]     A_reg_bank68_p0_rd_data;	// matmul/matmul-hw.mlir:12283:32
  wire [31:0]     A_reg_bank67_p0_rd_data;	// matmul/matmul-hw.mlir:12282:32
  wire [31:0]     A_reg_bank66_p0_rd_data;	// matmul/matmul-hw.mlir:12281:32
  wire [31:0]     A_reg_bank65_p0_rd_data;	// matmul/matmul-hw.mlir:12280:32
  wire [31:0]     A_reg_bank64_p0_rd_data;	// matmul/matmul-hw.mlir:12279:32
  wire [31:0]     A_reg_bank63_p0_rd_data;	// matmul/matmul-hw.mlir:12278:32
  wire [31:0]     A_reg_bank62_p0_rd_data;	// matmul/matmul-hw.mlir:12277:32
  wire [31:0]     A_reg_bank61_p0_rd_data;	// matmul/matmul-hw.mlir:12276:32
  wire [31:0]     A_reg_bank60_p0_rd_data;	// matmul/matmul-hw.mlir:12275:32
  wire [31:0]     A_reg_bank59_p0_rd_data;	// matmul/matmul-hw.mlir:12274:32
  wire [31:0]     A_reg_bank58_p0_rd_data;	// matmul/matmul-hw.mlir:12273:32
  wire [31:0]     A_reg_bank57_p0_rd_data;	// matmul/matmul-hw.mlir:12272:32
  wire [31:0]     A_reg_bank56_p0_rd_data;	// matmul/matmul-hw.mlir:12271:32
  wire [31:0]     A_reg_bank55_p0_rd_data;	// matmul/matmul-hw.mlir:12270:32
  wire [31:0]     A_reg_bank54_p0_rd_data;	// matmul/matmul-hw.mlir:12269:32
  wire [31:0]     A_reg_bank53_p0_rd_data;	// matmul/matmul-hw.mlir:12268:32
  wire [31:0]     A_reg_bank52_p0_rd_data;	// matmul/matmul-hw.mlir:12267:32
  wire [31:0]     A_reg_bank51_p0_rd_data;	// matmul/matmul-hw.mlir:12266:32
  wire [31:0]     A_reg_bank50_p0_rd_data;	// matmul/matmul-hw.mlir:12265:32
  wire [31:0]     A_reg_bank49_p0_rd_data;	// matmul/matmul-hw.mlir:12264:32
  wire [31:0]     A_reg_bank48_p0_rd_data;	// matmul/matmul-hw.mlir:12263:32
  wire [31:0]     A_reg_bank47_p0_rd_data;	// matmul/matmul-hw.mlir:12262:32
  wire [31:0]     A_reg_bank46_p0_rd_data;	// matmul/matmul-hw.mlir:12261:32
  wire [31:0]     A_reg_bank45_p0_rd_data;	// matmul/matmul-hw.mlir:12260:32
  wire [31:0]     A_reg_bank44_p0_rd_data;	// matmul/matmul-hw.mlir:12259:32
  wire [31:0]     A_reg_bank43_p0_rd_data;	// matmul/matmul-hw.mlir:12258:32
  wire [31:0]     A_reg_bank42_p0_rd_data;	// matmul/matmul-hw.mlir:12257:32
  wire [31:0]     A_reg_bank41_p0_rd_data;	// matmul/matmul-hw.mlir:12256:32
  wire [31:0]     A_reg_bank40_p0_rd_data;	// matmul/matmul-hw.mlir:12255:32
  wire [31:0]     A_reg_bank39_p0_rd_data;	// matmul/matmul-hw.mlir:12254:32
  wire [31:0]     A_reg_bank38_p0_rd_data;	// matmul/matmul-hw.mlir:12253:32
  wire [31:0]     A_reg_bank37_p0_rd_data;	// matmul/matmul-hw.mlir:12252:32
  wire [31:0]     A_reg_bank36_p0_rd_data;	// matmul/matmul-hw.mlir:12251:32
  wire [31:0]     A_reg_bank35_p0_rd_data;	// matmul/matmul-hw.mlir:12250:32
  wire [31:0]     A_reg_bank34_p0_rd_data;	// matmul/matmul-hw.mlir:12249:32
  wire [31:0]     A_reg_bank33_p0_rd_data;	// matmul/matmul-hw.mlir:12248:32
  wire [31:0]     A_reg_bank32_p0_rd_data;	// matmul/matmul-hw.mlir:12247:32
  wire [31:0]     A_reg_bank31_p0_rd_data;	// matmul/matmul-hw.mlir:12246:32
  wire [31:0]     A_reg_bank30_p0_rd_data;	// matmul/matmul-hw.mlir:12245:32
  wire [31:0]     A_reg_bank29_p0_rd_data;	// matmul/matmul-hw.mlir:12244:32
  wire [31:0]     A_reg_bank28_p0_rd_data;	// matmul/matmul-hw.mlir:12243:32
  wire [31:0]     A_reg_bank27_p0_rd_data;	// matmul/matmul-hw.mlir:12242:32
  wire [31:0]     A_reg_bank26_p0_rd_data;	// matmul/matmul-hw.mlir:12241:32
  wire [31:0]     A_reg_bank25_p0_rd_data;	// matmul/matmul-hw.mlir:12240:32
  wire [31:0]     A_reg_bank24_p0_rd_data;	// matmul/matmul-hw.mlir:12239:32
  wire [31:0]     A_reg_bank23_p0_rd_data;	// matmul/matmul-hw.mlir:12238:32
  wire [31:0]     A_reg_bank22_p0_rd_data;	// matmul/matmul-hw.mlir:12237:32
  wire [31:0]     A_reg_bank21_p0_rd_data;	// matmul/matmul-hw.mlir:12236:32
  wire [31:0]     A_reg_bank20_p0_rd_data;	// matmul/matmul-hw.mlir:12235:32
  wire [31:0]     A_reg_bank19_p0_rd_data;	// matmul/matmul-hw.mlir:12234:32
  wire [31:0]     A_reg_bank18_p0_rd_data;	// matmul/matmul-hw.mlir:12233:32
  wire [31:0]     A_reg_bank17_p0_rd_data;	// matmul/matmul-hw.mlir:12232:32
  wire [31:0]     A_reg_bank16_p0_rd_data;	// matmul/matmul-hw.mlir:12231:32
  wire [31:0]     A_reg_bank15_p0_rd_data;	// matmul/matmul-hw.mlir:12230:32
  wire [31:0]     A_reg_bank14_p0_rd_data;	// matmul/matmul-hw.mlir:12229:32
  wire [31:0]     A_reg_bank13_p0_rd_data;	// matmul/matmul-hw.mlir:12228:32
  wire [31:0]     A_reg_bank12_p0_rd_data;	// matmul/matmul-hw.mlir:12227:32
  wire [31:0]     A_reg_bank11_p0_rd_data;	// matmul/matmul-hw.mlir:12226:32
  wire [31:0]     A_reg_bank10_p0_rd_data;	// matmul/matmul-hw.mlir:12225:32
  wire [31:0]     A_reg_bank9_p0_rd_data;	// matmul/matmul-hw.mlir:12224:31
  wire [31:0]     A_reg_bank8_p0_rd_data;	// matmul/matmul-hw.mlir:12223:31
  wire [31:0]     A_reg_bank7_p0_rd_data;	// matmul/matmul-hw.mlir:12222:31
  wire [31:0]     A_reg_bank6_p0_rd_data;	// matmul/matmul-hw.mlir:12221:31
  wire [31:0]     A_reg_bank5_p0_rd_data;	// matmul/matmul-hw.mlir:12220:31
  wire [31:0]     A_reg_bank4_p0_rd_data;	// matmul/matmul-hw.mlir:12219:31
  wire [31:0]     A_reg_bank3_p0_rd_data;	// matmul/matmul-hw.mlir:12218:31
  wire [31:0]     A_reg_bank2_p0_rd_data;	// matmul/matmul-hw.mlir:12217:31
  wire [31:0]     A_reg_bank1_p0_rd_data;	// matmul/matmul-hw.mlir:12216:31
  wire [31:0]     A_reg_bank0_p0_rd_data;	// matmul/matmul-hw.mlir:12215:31
  wire            reg_1x1_r0_w1_inst3_p0_rd_data;	// matmul/matmul-hw.mlir:11178:39
  wire [5:0]      reg_1x6_r0_w1_inst3_p0_rd_data;	// matmul/matmul-hw.mlir:11167:39
  reg             _T_2710;	// matmul/matmul-hw.mlir:11144:12
  reg  [4:0]      _T_2716;	// matmul/matmul-hw.mlir:11183:12
  reg             _T_2719;	// matmul/matmul-hw.mlir:12475:12
  reg  [3:0]      i_k_next;	// matmul/matmul-hw.mlir:12493:17
  wire [3:0]      i_k_next_i_k_0;	// matmul/matmul-hw.mlir:12501:23
  reg  [1:0]      _T_2723;	// matmul/matmul-hw.mlir:12507:12
  reg  [1:0]      _T_2727;	// matmul/matmul-hw.mlir:12522:12
  reg  [3:0]      i_k_next_2732;	// matmul/matmul-hw.mlir:12539:22
  wire [3:0]      i_k_next_i_k_1;	// matmul/matmul-hw.mlir:12547:23
  reg  [2:0]      _T_2734;	// matmul/matmul-hw.mlir:12553:12
  reg  [2:0]      _T_2738;	// matmul/matmul-hw.mlir:12568:12
  reg  [3:0]      i_k_next_2743;	// matmul/matmul-hw.mlir:12585:22
  wire [3:0]      i_k_next_i_k_2;	// matmul/matmul-hw.mlir:12593:23
  reg  [3:0]      _T_2745;	// matmul/matmul-hw.mlir:12599:12
  reg  [3:0]      _T_2749;	// matmul/matmul-hw.mlir:12614:12
  reg  [3:0]      i_k_next_2754;	// matmul/matmul-hw.mlir:12631:22
  wire [3:0]      i_k_next_i_k_3;	// matmul/matmul-hw.mlir:12639:23
  reg  [4:0]      _T_2756;	// matmul/matmul-hw.mlir:12645:12
  reg  [4:0]      _T_2760;	// matmul/matmul-hw.mlir:12660:12
  reg  [3:0]      i_k_next_2765;	// matmul/matmul-hw.mlir:12677:22
  wire [3:0]      i_k_next_i_k_4;	// matmul/matmul-hw.mlir:12685:23
  reg  [5:0]      _T_2767;	// matmul/matmul-hw.mlir:12691:12
  reg  [5:0]      _T_2771;	// matmul/matmul-hw.mlir:12706:12
  reg  [3:0]      i_k_next_2776;	// matmul/matmul-hw.mlir:12723:22
  wire [3:0]      i_k_next_i_k_5;	// matmul/matmul-hw.mlir:12731:23
  reg  [6:0]      _T_2778;	// matmul/matmul-hw.mlir:12737:12
  reg  [6:0]      _T_2782;	// matmul/matmul-hw.mlir:12752:12
  reg  [3:0]      i_k_next_2787;	// matmul/matmul-hw.mlir:12769:22
  wire [3:0]      i_k_next_i_k_6;	// matmul/matmul-hw.mlir:12777:23
  reg  [7:0]      _T_2789;	// matmul/matmul-hw.mlir:12783:12
  reg  [7:0]      _T_2793;	// matmul/matmul-hw.mlir:12798:12
  reg  [3:0]      i_k_next_2798;	// matmul/matmul-hw.mlir:12815:22
  wire [3:0]      i_k_next_i_k_7;	// matmul/matmul-hw.mlir:12823:23
  reg  [8:0]      _T_2800;	// matmul/matmul-hw.mlir:12829:12
  reg  [8:0]      _T_2804;	// matmul/matmul-hw.mlir:12844:12
  reg  [3:0]      i_k_next_2809;	// matmul/matmul-hw.mlir:12861:22
  wire [3:0]      i_k_next_i_k_8;	// matmul/matmul-hw.mlir:12869:23
  reg  [9:0]      _T_2811;	// matmul/matmul-hw.mlir:12875:12
  reg  [9:0]      _T_2815;	// matmul/matmul-hw.mlir:12890:12
  reg  [3:0]      i_k_next_2820;	// matmul/matmul-hw.mlir:12907:22
  wire [3:0]      i_k_next_i_k_9;	// matmul/matmul-hw.mlir:12915:23
  reg  [10:0]     _T_2822;	// matmul/matmul-hw.mlir:12921:12
  reg  [10:0]     _T_2826;	// matmul/matmul-hw.mlir:12936:12
  reg  [3:0]      i_k_next_2831;	// matmul/matmul-hw.mlir:12953:22
  wire [3:0]      i_k_next_i_k_10;	// matmul/matmul-hw.mlir:12961:24
  reg  [11:0]     _T_2833;	// matmul/matmul-hw.mlir:12967:12
  reg  [11:0]     _T_2837;	// matmul/matmul-hw.mlir:12982:12
  reg  [3:0]      i_k_next_2842;	// matmul/matmul-hw.mlir:12999:22
  wire [3:0]      i_k_next_i_k_11;	// matmul/matmul-hw.mlir:13007:24
  reg  [12:0]     _T_2844;	// matmul/matmul-hw.mlir:13013:12
  reg  [12:0]     _T_2848;	// matmul/matmul-hw.mlir:13028:12
  reg  [3:0]      i_k_next_2853;	// matmul/matmul-hw.mlir:13045:22
  wire [3:0]      i_k_next_i_k_12;	// matmul/matmul-hw.mlir:13053:24
  reg  [13:0]     _T_2855;	// matmul/matmul-hw.mlir:13059:12
  reg  [13:0]     _T_2859;	// matmul/matmul-hw.mlir:13074:12
  reg  [3:0]      i_k_next_2864;	// matmul/matmul-hw.mlir:13091:22
  wire [3:0]      i_k_next_i_k_13;	// matmul/matmul-hw.mlir:13099:24
  reg  [14:0]     _T_2866;	// matmul/matmul-hw.mlir:13105:12
  reg  [14:0]     _T_2870;	// matmul/matmul-hw.mlir:13120:12
  reg  [3:0]      i_k_next_2875;	// matmul/matmul-hw.mlir:13137:22
  wire [3:0]      i_k_next_i_k_14;	// matmul/matmul-hw.mlir:13145:24
  reg  [15:0]     _T_2877;	// matmul/matmul-hw.mlir:13151:12
  reg  [15:0]     _T_2881;	// matmul/matmul-hw.mlir:13166:12
  reg  [3:0]      i_k_next_2886;	// matmul/matmul-hw.mlir:13183:22
  wire [3:0]      i_k_next_i_k_15;	// matmul/matmul-hw.mlir:13191:24
  reg  [16:0]     _T_2888;	// matmul/matmul-hw.mlir:13239:12
  reg  [17:0]     _T_2893;	// matmul/matmul-hw.mlir:13302:12
  reg  [18:0]     _T_2898;	// matmul/matmul-hw.mlir:13365:12
  reg  [19:0]     _T_2903;	// matmul/matmul-hw.mlir:13428:12
  reg  [20:0]     _T_2908;	// matmul/matmul-hw.mlir:13491:12
  reg  [21:0]     _T_2913;	// matmul/matmul-hw.mlir:13554:12
  reg  [22:0]     _T_2918;	// matmul/matmul-hw.mlir:13617:12
  reg  [23:0]     _T_2923;	// matmul/matmul-hw.mlir:13680:13
  reg  [24:0]     _T_2928;	// matmul/matmul-hw.mlir:13743:13
  reg  [25:0]     _T_2933;	// matmul/matmul-hw.mlir:13806:13
  reg  [26:0]     _T_2938;	// matmul/matmul-hw.mlir:13869:13
  reg  [27:0]     _T_2943;	// matmul/matmul-hw.mlir:13932:13
  reg  [28:0]     _T_2948;	// matmul/matmul-hw.mlir:13995:13
  reg  [29:0]     _T_2953;	// matmul/matmul-hw.mlir:14058:13
  reg  [30:0]     _T_2958;	// matmul/matmul-hw.mlir:14121:13
  wire [31:0]     a_i_k_0_i_j_0;	// matmul/matmul-hw.mlir:14230:22
  wire [31:0]     b_i_k_0_i_j_0;	// matmul/matmul-hw.mlir:14233:22
  wire [31:0]     c_prev_i_k_0_i_j_0;	// matmul/matmul-hw.mlir:14236:27
  wire            tk_i_k_0_i_j_0;	// matmul/matmul-hw.mlir:14239:23
  wire [31:0]     c_i_k_0_i_j_0;	// matmul/matmul-hw.mlir:14243:22
  wire [31:0]     a_i_k_1_i_j_0;	// matmul/matmul-hw.mlir:14252:22
  wire [31:0]     b_i_k_1_i_j_0;	// matmul/matmul-hw.mlir:14255:22
  wire [31:0]     c_prev_i_k_1_i_j_0;	// matmul/matmul-hw.mlir:14258:27
  wire            tk_i_k_1_i_j_0;	// matmul/matmul-hw.mlir:14261:23
  wire [31:0]     c_i_k_1_i_j_0;	// matmul/matmul-hw.mlir:14265:22
  wire [31:0]     a_i_k_2_i_j_0;	// matmul/matmul-hw.mlir:14274:22
  wire [31:0]     b_i_k_2_i_j_0;	// matmul/matmul-hw.mlir:14277:22
  wire [31:0]     c_prev_i_k_2_i_j_0;	// matmul/matmul-hw.mlir:14280:27
  wire            tk_i_k_2_i_j_0;	// matmul/matmul-hw.mlir:14283:23
  wire [31:0]     c_i_k_2_i_j_0;	// matmul/matmul-hw.mlir:14287:22
  wire [31:0]     a_i_k_3_i_j_0;	// matmul/matmul-hw.mlir:14296:22
  wire [31:0]     b_i_k_3_i_j_0;	// matmul/matmul-hw.mlir:14299:22
  wire [31:0]     c_prev_i_k_3_i_j_0;	// matmul/matmul-hw.mlir:14302:27
  wire            tk_i_k_3_i_j_0;	// matmul/matmul-hw.mlir:14305:23
  wire [31:0]     c_i_k_3_i_j_0;	// matmul/matmul-hw.mlir:14309:22
  wire [31:0]     a_i_k_4_i_j_0;	// matmul/matmul-hw.mlir:14318:22
  wire [31:0]     b_i_k_4_i_j_0;	// matmul/matmul-hw.mlir:14321:22
  wire [31:0]     c_prev_i_k_4_i_j_0;	// matmul/matmul-hw.mlir:14324:27
  wire            tk_i_k_4_i_j_0;	// matmul/matmul-hw.mlir:14327:23
  wire [31:0]     c_i_k_4_i_j_0;	// matmul/matmul-hw.mlir:14331:22
  wire [31:0]     a_i_k_5_i_j_0;	// matmul/matmul-hw.mlir:14340:22
  wire [31:0]     b_i_k_5_i_j_0;	// matmul/matmul-hw.mlir:14343:22
  wire [31:0]     c_prev_i_k_5_i_j_0;	// matmul/matmul-hw.mlir:14346:27
  wire            tk_i_k_5_i_j_0;	// matmul/matmul-hw.mlir:14349:23
  wire [31:0]     c_i_k_5_i_j_0;	// matmul/matmul-hw.mlir:14353:22
  wire [31:0]     a_i_k_6_i_j_0;	// matmul/matmul-hw.mlir:14362:22
  wire [31:0]     b_i_k_6_i_j_0;	// matmul/matmul-hw.mlir:14365:22
  wire [31:0]     c_prev_i_k_6_i_j_0;	// matmul/matmul-hw.mlir:14368:27
  wire            tk_i_k_6_i_j_0;	// matmul/matmul-hw.mlir:14371:23
  wire [31:0]     c_i_k_6_i_j_0;	// matmul/matmul-hw.mlir:14375:22
  wire [31:0]     a_i_k_7_i_j_0;	// matmul/matmul-hw.mlir:14384:22
  wire [31:0]     b_i_k_7_i_j_0;	// matmul/matmul-hw.mlir:14387:22
  wire [31:0]     c_prev_i_k_7_i_j_0;	// matmul/matmul-hw.mlir:14390:27
  wire            tk_i_k_7_i_j_0;	// matmul/matmul-hw.mlir:14393:23
  wire [31:0]     c_i_k_7_i_j_0;	// matmul/matmul-hw.mlir:14397:22
  wire [31:0]     a_i_k_8_i_j_0;	// matmul/matmul-hw.mlir:14406:22
  wire [31:0]     b_i_k_8_i_j_0;	// matmul/matmul-hw.mlir:14409:22
  wire [31:0]     c_prev_i_k_8_i_j_0;	// matmul/matmul-hw.mlir:14412:27
  wire            tk_i_k_8_i_j_0;	// matmul/matmul-hw.mlir:14415:23
  wire [31:0]     c_i_k_8_i_j_0;	// matmul/matmul-hw.mlir:14419:22
  wire [31:0]     a_i_k_9_i_j_0;	// matmul/matmul-hw.mlir:14428:22
  wire [31:0]     b_i_k_9_i_j_0;	// matmul/matmul-hw.mlir:14431:22
  wire [31:0]     c_prev_i_k_9_i_j_0;	// matmul/matmul-hw.mlir:14434:27
  wire            tk_i_k_9_i_j_0;	// matmul/matmul-hw.mlir:14437:23
  wire [31:0]     c_i_k_9_i_j_0;	// matmul/matmul-hw.mlir:14441:22
  wire [31:0]     a_i_k_10_i_j_0;	// matmul/matmul-hw.mlir:14450:23
  wire [31:0]     b_i_k_10_i_j_0;	// matmul/matmul-hw.mlir:14453:23
  wire [31:0]     c_prev_i_k_10_i_j_0;	// matmul/matmul-hw.mlir:14456:28
  wire            tk_i_k_10_i_j_0;	// matmul/matmul-hw.mlir:14459:24
  wire [31:0]     c_i_k_10_i_j_0;	// matmul/matmul-hw.mlir:14463:23
  wire [31:0]     a_i_k_11_i_j_0;	// matmul/matmul-hw.mlir:14472:23
  wire [31:0]     b_i_k_11_i_j_0;	// matmul/matmul-hw.mlir:14475:23
  wire [31:0]     c_prev_i_k_11_i_j_0;	// matmul/matmul-hw.mlir:14478:28
  wire            tk_i_k_11_i_j_0;	// matmul/matmul-hw.mlir:14481:24
  wire [31:0]     c_i_k_11_i_j_0;	// matmul/matmul-hw.mlir:14485:23
  wire [31:0]     a_i_k_12_i_j_0;	// matmul/matmul-hw.mlir:14494:23
  wire [31:0]     b_i_k_12_i_j_0;	// matmul/matmul-hw.mlir:14497:23
  wire [31:0]     c_prev_i_k_12_i_j_0;	// matmul/matmul-hw.mlir:14500:28
  wire            tk_i_k_12_i_j_0;	// matmul/matmul-hw.mlir:14503:24
  wire [31:0]     c_i_k_12_i_j_0;	// matmul/matmul-hw.mlir:14507:23
  wire [31:0]     a_i_k_13_i_j_0;	// matmul/matmul-hw.mlir:14516:23
  wire [31:0]     b_i_k_13_i_j_0;	// matmul/matmul-hw.mlir:14519:23
  wire [31:0]     c_prev_i_k_13_i_j_0;	// matmul/matmul-hw.mlir:14522:28
  wire            tk_i_k_13_i_j_0;	// matmul/matmul-hw.mlir:14525:24
  wire [31:0]     c_i_k_13_i_j_0;	// matmul/matmul-hw.mlir:14529:23
  wire [31:0]     a_i_k_14_i_j_0;	// matmul/matmul-hw.mlir:14538:23
  wire [31:0]     b_i_k_14_i_j_0;	// matmul/matmul-hw.mlir:14541:23
  wire [31:0]     c_prev_i_k_14_i_j_0;	// matmul/matmul-hw.mlir:14544:28
  wire            tk_i_k_14_i_j_0;	// matmul/matmul-hw.mlir:14547:24
  wire [31:0]     c_i_k_14_i_j_0;	// matmul/matmul-hw.mlir:14551:23
  wire [31:0]     a_i_k_15_i_j_0;	// matmul/matmul-hw.mlir:14560:23
  wire [31:0]     b_i_k_15_i_j_0;	// matmul/matmul-hw.mlir:14563:23
  wire [31:0]     c_prev_i_k_15_i_j_0;	// matmul/matmul-hw.mlir:14566:28
  wire            tk_i_k_15_i_j_0;	// matmul/matmul-hw.mlir:14569:24
  wire [31:0]     c_i_k_15_i_j_0;	// matmul/matmul-hw.mlir:14573:23
  reg  [3:0][3:0] i_delayed;	// matmul/matmul-hw.mlir:14579:18
  reg  [3:0]      i_j_next;	// matmul/matmul-hw.mlir:14598:17
  wire [31:0]     a_i_k_0_i_j_1;	// matmul/matmul-hw.mlir:14697:22
  wire [31:0]     b_i_k_0_i_j_1;	// matmul/matmul-hw.mlir:14700:22
  wire [31:0]     c_prev_i_k_0_i_j_1;	// matmul/matmul-hw.mlir:14703:27
  wire            tk_i_k_0_i_j_1;	// matmul/matmul-hw.mlir:14706:23
  wire [31:0]     c_i_k_0_i_j_1;	// matmul/matmul-hw.mlir:14710:22
  reg  [3:0]      i_k_next_3001;	// matmul/matmul-hw.mlir:14715:22
  wire [31:0]     a_i_k_1_i_j_1;	// matmul/matmul-hw.mlir:14727:22
  wire [31:0]     b_i_k_1_i_j_1;	// matmul/matmul-hw.mlir:14730:22
  wire [31:0]     c_prev_i_k_1_i_j_1;	// matmul/matmul-hw.mlir:14733:27
  wire            tk_i_k_1_i_j_1;	// matmul/matmul-hw.mlir:14736:23
  wire [31:0]     c_i_k_1_i_j_1;	// matmul/matmul-hw.mlir:14740:22
  reg  [3:0]      i_k_next_3004;	// matmul/matmul-hw.mlir:14745:22
  wire [31:0]     a_i_k_2_i_j_1;	// matmul/matmul-hw.mlir:14757:22
  wire [31:0]     b_i_k_2_i_j_1;	// matmul/matmul-hw.mlir:14760:22
  wire [31:0]     c_prev_i_k_2_i_j_1;	// matmul/matmul-hw.mlir:14763:27
  wire            tk_i_k_2_i_j_1;	// matmul/matmul-hw.mlir:14766:23
  wire [31:0]     c_i_k_2_i_j_1;	// matmul/matmul-hw.mlir:14770:22
  reg  [3:0]      i_k_next_3007;	// matmul/matmul-hw.mlir:14775:22
  wire [31:0]     a_i_k_3_i_j_1;	// matmul/matmul-hw.mlir:14787:22
  wire [31:0]     b_i_k_3_i_j_1;	// matmul/matmul-hw.mlir:14790:22
  wire [31:0]     c_prev_i_k_3_i_j_1;	// matmul/matmul-hw.mlir:14793:27
  wire            tk_i_k_3_i_j_1;	// matmul/matmul-hw.mlir:14796:23
  wire [31:0]     c_i_k_3_i_j_1;	// matmul/matmul-hw.mlir:14800:22
  reg  [3:0]      i_k_next_3010;	// matmul/matmul-hw.mlir:14805:22
  wire [31:0]     a_i_k_4_i_j_1;	// matmul/matmul-hw.mlir:14817:22
  wire [31:0]     b_i_k_4_i_j_1;	// matmul/matmul-hw.mlir:14820:22
  wire [31:0]     c_prev_i_k_4_i_j_1;	// matmul/matmul-hw.mlir:14823:27
  wire            tk_i_k_4_i_j_1;	// matmul/matmul-hw.mlir:14826:23
  wire [31:0]     c_i_k_4_i_j_1;	// matmul/matmul-hw.mlir:14830:22
  reg  [3:0]      i_k_next_3013;	// matmul/matmul-hw.mlir:14835:22
  wire [31:0]     a_i_k_5_i_j_1;	// matmul/matmul-hw.mlir:14847:22
  wire [31:0]     b_i_k_5_i_j_1;	// matmul/matmul-hw.mlir:14850:22
  wire [31:0]     c_prev_i_k_5_i_j_1;	// matmul/matmul-hw.mlir:14853:27
  wire            tk_i_k_5_i_j_1;	// matmul/matmul-hw.mlir:14856:23
  wire [31:0]     c_i_k_5_i_j_1;	// matmul/matmul-hw.mlir:14860:22
  reg  [3:0]      i_k_next_3016;	// matmul/matmul-hw.mlir:14865:22
  wire [31:0]     a_i_k_6_i_j_1;	// matmul/matmul-hw.mlir:14877:22
  wire [31:0]     b_i_k_6_i_j_1;	// matmul/matmul-hw.mlir:14880:22
  wire [31:0]     c_prev_i_k_6_i_j_1;	// matmul/matmul-hw.mlir:14883:27
  wire            tk_i_k_6_i_j_1;	// matmul/matmul-hw.mlir:14886:23
  wire [31:0]     c_i_k_6_i_j_1;	// matmul/matmul-hw.mlir:14890:22
  reg  [3:0]      i_k_next_3019;	// matmul/matmul-hw.mlir:14895:22
  wire [31:0]     a_i_k_7_i_j_1;	// matmul/matmul-hw.mlir:14907:22
  wire [31:0]     b_i_k_7_i_j_1;	// matmul/matmul-hw.mlir:14910:22
  wire [31:0]     c_prev_i_k_7_i_j_1;	// matmul/matmul-hw.mlir:14913:27
  wire            tk_i_k_7_i_j_1;	// matmul/matmul-hw.mlir:14916:23
  wire [31:0]     c_i_k_7_i_j_1;	// matmul/matmul-hw.mlir:14920:22
  reg  [3:0]      i_k_next_3022;	// matmul/matmul-hw.mlir:14925:22
  wire [31:0]     a_i_k_8_i_j_1;	// matmul/matmul-hw.mlir:14937:22
  wire [31:0]     b_i_k_8_i_j_1;	// matmul/matmul-hw.mlir:14940:22
  wire [31:0]     c_prev_i_k_8_i_j_1;	// matmul/matmul-hw.mlir:14943:27
  wire            tk_i_k_8_i_j_1;	// matmul/matmul-hw.mlir:14946:23
  wire [31:0]     c_i_k_8_i_j_1;	// matmul/matmul-hw.mlir:14950:22
  reg  [3:0]      i_k_next_3025;	// matmul/matmul-hw.mlir:14955:22
  wire [31:0]     a_i_k_9_i_j_1;	// matmul/matmul-hw.mlir:14967:22
  wire [31:0]     b_i_k_9_i_j_1;	// matmul/matmul-hw.mlir:14970:22
  wire [31:0]     c_prev_i_k_9_i_j_1;	// matmul/matmul-hw.mlir:14973:27
  wire            tk_i_k_9_i_j_1;	// matmul/matmul-hw.mlir:14976:23
  wire [31:0]     c_i_k_9_i_j_1;	// matmul/matmul-hw.mlir:14980:22
  reg  [3:0]      i_k_next_3028;	// matmul/matmul-hw.mlir:14985:22
  wire [31:0]     a_i_k_10_i_j_1;	// matmul/matmul-hw.mlir:14997:23
  wire [31:0]     b_i_k_10_i_j_1;	// matmul/matmul-hw.mlir:15000:23
  wire [31:0]     c_prev_i_k_10_i_j_1;	// matmul/matmul-hw.mlir:15003:28
  wire            tk_i_k_10_i_j_1;	// matmul/matmul-hw.mlir:15006:24
  wire [31:0]     c_i_k_10_i_j_1;	// matmul/matmul-hw.mlir:15010:23
  reg  [3:0]      i_k_next_3031;	// matmul/matmul-hw.mlir:15015:22
  wire [31:0]     a_i_k_11_i_j_1;	// matmul/matmul-hw.mlir:15027:23
  wire [31:0]     b_i_k_11_i_j_1;	// matmul/matmul-hw.mlir:15030:23
  wire [31:0]     c_prev_i_k_11_i_j_1;	// matmul/matmul-hw.mlir:15033:28
  wire            tk_i_k_11_i_j_1;	// matmul/matmul-hw.mlir:15036:24
  wire [31:0]     c_i_k_11_i_j_1;	// matmul/matmul-hw.mlir:15040:23
  reg  [3:0]      i_k_next_3034;	// matmul/matmul-hw.mlir:15045:22
  wire [31:0]     a_i_k_12_i_j_1;	// matmul/matmul-hw.mlir:15057:23
  wire [31:0]     b_i_k_12_i_j_1;	// matmul/matmul-hw.mlir:15060:23
  wire [31:0]     c_prev_i_k_12_i_j_1;	// matmul/matmul-hw.mlir:15063:28
  wire            tk_i_k_12_i_j_1;	// matmul/matmul-hw.mlir:15066:24
  wire [31:0]     c_i_k_12_i_j_1;	// matmul/matmul-hw.mlir:15070:23
  reg  [3:0]      i_k_next_3037;	// matmul/matmul-hw.mlir:15075:22
  wire [31:0]     a_i_k_13_i_j_1;	// matmul/matmul-hw.mlir:15087:23
  wire [31:0]     b_i_k_13_i_j_1;	// matmul/matmul-hw.mlir:15090:23
  wire [31:0]     c_prev_i_k_13_i_j_1;	// matmul/matmul-hw.mlir:15093:28
  wire            tk_i_k_13_i_j_1;	// matmul/matmul-hw.mlir:15096:24
  wire [31:0]     c_i_k_13_i_j_1;	// matmul/matmul-hw.mlir:15100:23
  reg  [3:0]      i_k_next_3040;	// matmul/matmul-hw.mlir:15105:22
  wire [31:0]     a_i_k_14_i_j_1;	// matmul/matmul-hw.mlir:15117:23
  wire [31:0]     b_i_k_14_i_j_1;	// matmul/matmul-hw.mlir:15120:23
  wire [31:0]     c_prev_i_k_14_i_j_1;	// matmul/matmul-hw.mlir:15123:28
  wire            tk_i_k_14_i_j_1;	// matmul/matmul-hw.mlir:15126:24
  wire [31:0]     c_i_k_14_i_j_1;	// matmul/matmul-hw.mlir:15130:23
  reg  [3:0]      i_k_next_3043;	// matmul/matmul-hw.mlir:15135:22
  wire [31:0]     a_i_k_15_i_j_1;	// matmul/matmul-hw.mlir:15147:23
  wire [31:0]     b_i_k_15_i_j_1;	// matmul/matmul-hw.mlir:15150:23
  wire [31:0]     c_prev_i_k_15_i_j_1;	// matmul/matmul-hw.mlir:15153:28
  wire            tk_i_k_15_i_j_1;	// matmul/matmul-hw.mlir:15156:24
  wire [31:0]     c_i_k_15_i_j_1;	// matmul/matmul-hw.mlir:15160:23
  reg  [3:0]      i_k_next_3046;	// matmul/matmul-hw.mlir:15165:22
  reg  [3:0][3:0] i_delayed_3048;	// matmul/matmul-hw.mlir:15174:23
  reg  [3:0]      i_j_next_3052;	// matmul/matmul-hw.mlir:15193:22
  wire [31:0]     a_i_k_0_i_j_2;	// matmul/matmul-hw.mlir:15292:22
  wire [31:0]     b_i_k_0_i_j_2;	// matmul/matmul-hw.mlir:15295:22
  wire [31:0]     c_prev_i_k_0_i_j_2;	// matmul/matmul-hw.mlir:15298:27
  wire            tk_i_k_0_i_j_2;	// matmul/matmul-hw.mlir:15301:23
  wire [31:0]     c_i_k_0_i_j_2;	// matmul/matmul-hw.mlir:15305:22
  reg  [3:0]      i_k_next_3072;	// matmul/matmul-hw.mlir:15310:22
  wire [31:0]     a_i_k_1_i_j_2;	// matmul/matmul-hw.mlir:15322:22
  wire [31:0]     b_i_k_1_i_j_2;	// matmul/matmul-hw.mlir:15325:22
  wire [31:0]     c_prev_i_k_1_i_j_2;	// matmul/matmul-hw.mlir:15328:27
  wire            tk_i_k_1_i_j_2;	// matmul/matmul-hw.mlir:15331:23
  wire [31:0]     c_i_k_1_i_j_2;	// matmul/matmul-hw.mlir:15335:22
  reg  [3:0]      i_k_next_3075;	// matmul/matmul-hw.mlir:15340:22
  wire [31:0]     a_i_k_2_i_j_2;	// matmul/matmul-hw.mlir:15352:22
  wire [31:0]     b_i_k_2_i_j_2;	// matmul/matmul-hw.mlir:15355:22
  wire [31:0]     c_prev_i_k_2_i_j_2;	// matmul/matmul-hw.mlir:15358:27
  wire            tk_i_k_2_i_j_2;	// matmul/matmul-hw.mlir:15361:23
  wire [31:0]     c_i_k_2_i_j_2;	// matmul/matmul-hw.mlir:15365:22
  reg  [3:0]      i_k_next_3078;	// matmul/matmul-hw.mlir:15370:22
  wire [31:0]     a_i_k_3_i_j_2;	// matmul/matmul-hw.mlir:15382:22
  wire [31:0]     b_i_k_3_i_j_2;	// matmul/matmul-hw.mlir:15385:22
  wire [31:0]     c_prev_i_k_3_i_j_2;	// matmul/matmul-hw.mlir:15388:27
  wire            tk_i_k_3_i_j_2;	// matmul/matmul-hw.mlir:15391:23
  wire [31:0]     c_i_k_3_i_j_2;	// matmul/matmul-hw.mlir:15395:22
  reg  [3:0]      i_k_next_3081;	// matmul/matmul-hw.mlir:15400:22
  wire [31:0]     a_i_k_4_i_j_2;	// matmul/matmul-hw.mlir:15412:22
  wire [31:0]     b_i_k_4_i_j_2;	// matmul/matmul-hw.mlir:15415:22
  wire [31:0]     c_prev_i_k_4_i_j_2;	// matmul/matmul-hw.mlir:15418:27
  wire            tk_i_k_4_i_j_2;	// matmul/matmul-hw.mlir:15421:23
  wire [31:0]     c_i_k_4_i_j_2;	// matmul/matmul-hw.mlir:15425:22
  reg  [3:0]      i_k_next_3084;	// matmul/matmul-hw.mlir:15430:22
  wire [31:0]     a_i_k_5_i_j_2;	// matmul/matmul-hw.mlir:15442:22
  wire [31:0]     b_i_k_5_i_j_2;	// matmul/matmul-hw.mlir:15445:22
  wire [31:0]     c_prev_i_k_5_i_j_2;	// matmul/matmul-hw.mlir:15448:27
  wire            tk_i_k_5_i_j_2;	// matmul/matmul-hw.mlir:15451:23
  wire [31:0]     c_i_k_5_i_j_2;	// matmul/matmul-hw.mlir:15455:22
  reg  [3:0]      i_k_next_3087;	// matmul/matmul-hw.mlir:15460:22
  wire [31:0]     a_i_k_6_i_j_2;	// matmul/matmul-hw.mlir:15472:22
  wire [31:0]     b_i_k_6_i_j_2;	// matmul/matmul-hw.mlir:15475:22
  wire [31:0]     c_prev_i_k_6_i_j_2;	// matmul/matmul-hw.mlir:15478:27
  wire            tk_i_k_6_i_j_2;	// matmul/matmul-hw.mlir:15481:23
  wire [31:0]     c_i_k_6_i_j_2;	// matmul/matmul-hw.mlir:15485:22
  reg  [3:0]      i_k_next_3090;	// matmul/matmul-hw.mlir:15490:22
  wire [31:0]     a_i_k_7_i_j_2;	// matmul/matmul-hw.mlir:15502:22
  wire [31:0]     b_i_k_7_i_j_2;	// matmul/matmul-hw.mlir:15505:22
  wire [31:0]     c_prev_i_k_7_i_j_2;	// matmul/matmul-hw.mlir:15508:27
  wire            tk_i_k_7_i_j_2;	// matmul/matmul-hw.mlir:15511:23
  wire [31:0]     c_i_k_7_i_j_2;	// matmul/matmul-hw.mlir:15515:22
  reg  [3:0]      i_k_next_3093;	// matmul/matmul-hw.mlir:15520:22
  wire [31:0]     a_i_k_8_i_j_2;	// matmul/matmul-hw.mlir:15532:22
  wire [31:0]     b_i_k_8_i_j_2;	// matmul/matmul-hw.mlir:15535:22
  wire [31:0]     c_prev_i_k_8_i_j_2;	// matmul/matmul-hw.mlir:15538:27
  wire            tk_i_k_8_i_j_2;	// matmul/matmul-hw.mlir:15541:23
  wire [31:0]     c_i_k_8_i_j_2;	// matmul/matmul-hw.mlir:15545:22
  reg  [3:0]      i_k_next_3096;	// matmul/matmul-hw.mlir:15550:22
  wire [31:0]     a_i_k_9_i_j_2;	// matmul/matmul-hw.mlir:15562:22
  wire [31:0]     b_i_k_9_i_j_2;	// matmul/matmul-hw.mlir:15565:22
  wire [31:0]     c_prev_i_k_9_i_j_2;	// matmul/matmul-hw.mlir:15568:27
  wire            tk_i_k_9_i_j_2;	// matmul/matmul-hw.mlir:15571:23
  wire [31:0]     c_i_k_9_i_j_2;	// matmul/matmul-hw.mlir:15575:22
  reg  [3:0]      i_k_next_3099;	// matmul/matmul-hw.mlir:15580:22
  wire [31:0]     a_i_k_10_i_j_2;	// matmul/matmul-hw.mlir:15592:23
  wire [31:0]     b_i_k_10_i_j_2;	// matmul/matmul-hw.mlir:15595:23
  wire [31:0]     c_prev_i_k_10_i_j_2;	// matmul/matmul-hw.mlir:15598:28
  wire            tk_i_k_10_i_j_2;	// matmul/matmul-hw.mlir:15601:24
  wire [31:0]     c_i_k_10_i_j_2;	// matmul/matmul-hw.mlir:15605:23
  reg  [3:0]      i_k_next_3102;	// matmul/matmul-hw.mlir:15610:22
  wire [31:0]     a_i_k_11_i_j_2;	// matmul/matmul-hw.mlir:15622:23
  wire [31:0]     b_i_k_11_i_j_2;	// matmul/matmul-hw.mlir:15625:23
  wire [31:0]     c_prev_i_k_11_i_j_2;	// matmul/matmul-hw.mlir:15628:28
  wire            tk_i_k_11_i_j_2;	// matmul/matmul-hw.mlir:15631:24
  wire [31:0]     c_i_k_11_i_j_2;	// matmul/matmul-hw.mlir:15635:23
  reg  [3:0]      i_k_next_3105;	// matmul/matmul-hw.mlir:15640:22
  wire [31:0]     a_i_k_12_i_j_2;	// matmul/matmul-hw.mlir:15652:23
  wire [31:0]     b_i_k_12_i_j_2;	// matmul/matmul-hw.mlir:15655:23
  wire [31:0]     c_prev_i_k_12_i_j_2;	// matmul/matmul-hw.mlir:15658:28
  wire            tk_i_k_12_i_j_2;	// matmul/matmul-hw.mlir:15661:24
  wire [31:0]     c_i_k_12_i_j_2;	// matmul/matmul-hw.mlir:15665:23
  reg  [3:0]      i_k_next_3108;	// matmul/matmul-hw.mlir:15670:22
  wire [31:0]     a_i_k_13_i_j_2;	// matmul/matmul-hw.mlir:15682:23
  wire [31:0]     b_i_k_13_i_j_2;	// matmul/matmul-hw.mlir:15685:23
  wire [31:0]     c_prev_i_k_13_i_j_2;	// matmul/matmul-hw.mlir:15688:28
  wire            tk_i_k_13_i_j_2;	// matmul/matmul-hw.mlir:15691:24
  wire [31:0]     c_i_k_13_i_j_2;	// matmul/matmul-hw.mlir:15695:23
  reg  [3:0]      i_k_next_3111;	// matmul/matmul-hw.mlir:15700:22
  wire [31:0]     a_i_k_14_i_j_2;	// matmul/matmul-hw.mlir:15712:23
  wire [31:0]     b_i_k_14_i_j_2;	// matmul/matmul-hw.mlir:15715:23
  wire [31:0]     c_prev_i_k_14_i_j_2;	// matmul/matmul-hw.mlir:15718:28
  wire            tk_i_k_14_i_j_2;	// matmul/matmul-hw.mlir:15721:24
  wire [31:0]     c_i_k_14_i_j_2;	// matmul/matmul-hw.mlir:15725:23
  reg  [3:0]      i_k_next_3114;	// matmul/matmul-hw.mlir:15730:22
  wire [31:0]     a_i_k_15_i_j_2;	// matmul/matmul-hw.mlir:15742:23
  wire [31:0]     b_i_k_15_i_j_2;	// matmul/matmul-hw.mlir:15745:23
  wire [31:0]     c_prev_i_k_15_i_j_2;	// matmul/matmul-hw.mlir:15748:28
  wire            tk_i_k_15_i_j_2;	// matmul/matmul-hw.mlir:15751:24
  wire [31:0]     c_i_k_15_i_j_2;	// matmul/matmul-hw.mlir:15755:23
  reg  [3:0]      i_k_next_3117;	// matmul/matmul-hw.mlir:15760:22
  reg  [3:0][3:0] i_delayed_3119;	// matmul/matmul-hw.mlir:15769:23
  reg  [3:0]      i_j_next_3123;	// matmul/matmul-hw.mlir:15788:22
  wire [31:0]     a_i_k_0_i_j_3;	// matmul/matmul-hw.mlir:15887:22
  wire [31:0]     b_i_k_0_i_j_3;	// matmul/matmul-hw.mlir:15890:22
  wire [31:0]     c_prev_i_k_0_i_j_3;	// matmul/matmul-hw.mlir:15893:27
  wire            tk_i_k_0_i_j_3;	// matmul/matmul-hw.mlir:15896:23
  wire [31:0]     c_i_k_0_i_j_3;	// matmul/matmul-hw.mlir:15900:22
  reg  [3:0]      i_k_next_3143;	// matmul/matmul-hw.mlir:15905:22
  wire [31:0]     a_i_k_1_i_j_3;	// matmul/matmul-hw.mlir:15917:22
  wire [31:0]     b_i_k_1_i_j_3;	// matmul/matmul-hw.mlir:15920:22
  wire [31:0]     c_prev_i_k_1_i_j_3;	// matmul/matmul-hw.mlir:15923:27
  wire            tk_i_k_1_i_j_3;	// matmul/matmul-hw.mlir:15926:23
  wire [31:0]     c_i_k_1_i_j_3;	// matmul/matmul-hw.mlir:15930:22
  reg  [3:0]      i_k_next_3146;	// matmul/matmul-hw.mlir:15935:22
  wire [31:0]     a_i_k_2_i_j_3;	// matmul/matmul-hw.mlir:15947:22
  wire [31:0]     b_i_k_2_i_j_3;	// matmul/matmul-hw.mlir:15950:22
  wire [31:0]     c_prev_i_k_2_i_j_3;	// matmul/matmul-hw.mlir:15953:27
  wire            tk_i_k_2_i_j_3;	// matmul/matmul-hw.mlir:15956:23
  wire [31:0]     c_i_k_2_i_j_3;	// matmul/matmul-hw.mlir:15960:22
  reg  [3:0]      i_k_next_3149;	// matmul/matmul-hw.mlir:15965:22
  wire [31:0]     a_i_k_3_i_j_3;	// matmul/matmul-hw.mlir:15977:22
  wire [31:0]     b_i_k_3_i_j_3;	// matmul/matmul-hw.mlir:15980:22
  wire [31:0]     c_prev_i_k_3_i_j_3;	// matmul/matmul-hw.mlir:15983:27
  wire            tk_i_k_3_i_j_3;	// matmul/matmul-hw.mlir:15986:23
  wire [31:0]     c_i_k_3_i_j_3;	// matmul/matmul-hw.mlir:15990:22
  reg  [3:0]      i_k_next_3152;	// matmul/matmul-hw.mlir:15995:22
  wire [31:0]     a_i_k_4_i_j_3;	// matmul/matmul-hw.mlir:16007:22
  wire [31:0]     b_i_k_4_i_j_3;	// matmul/matmul-hw.mlir:16010:22
  wire [31:0]     c_prev_i_k_4_i_j_3;	// matmul/matmul-hw.mlir:16013:27
  wire            tk_i_k_4_i_j_3;	// matmul/matmul-hw.mlir:16016:23
  wire [31:0]     c_i_k_4_i_j_3;	// matmul/matmul-hw.mlir:16020:22
  reg  [3:0]      i_k_next_3155;	// matmul/matmul-hw.mlir:16025:22
  wire [31:0]     a_i_k_5_i_j_3;	// matmul/matmul-hw.mlir:16037:22
  wire [31:0]     b_i_k_5_i_j_3;	// matmul/matmul-hw.mlir:16040:22
  wire [31:0]     c_prev_i_k_5_i_j_3;	// matmul/matmul-hw.mlir:16043:27
  wire            tk_i_k_5_i_j_3;	// matmul/matmul-hw.mlir:16046:23
  wire [31:0]     c_i_k_5_i_j_3;	// matmul/matmul-hw.mlir:16050:22
  reg  [3:0]      i_k_next_3158;	// matmul/matmul-hw.mlir:16055:22
  wire [31:0]     a_i_k_6_i_j_3;	// matmul/matmul-hw.mlir:16067:22
  wire [31:0]     b_i_k_6_i_j_3;	// matmul/matmul-hw.mlir:16070:22
  wire [31:0]     c_prev_i_k_6_i_j_3;	// matmul/matmul-hw.mlir:16073:27
  wire            tk_i_k_6_i_j_3;	// matmul/matmul-hw.mlir:16076:23
  wire [31:0]     c_i_k_6_i_j_3;	// matmul/matmul-hw.mlir:16080:22
  reg  [3:0]      i_k_next_3161;	// matmul/matmul-hw.mlir:16085:22
  wire [31:0]     a_i_k_7_i_j_3;	// matmul/matmul-hw.mlir:16097:22
  wire [31:0]     b_i_k_7_i_j_3;	// matmul/matmul-hw.mlir:16100:22
  wire [31:0]     c_prev_i_k_7_i_j_3;	// matmul/matmul-hw.mlir:16103:27
  wire            tk_i_k_7_i_j_3;	// matmul/matmul-hw.mlir:16106:23
  wire [31:0]     c_i_k_7_i_j_3;	// matmul/matmul-hw.mlir:16110:22
  reg  [3:0]      i_k_next_3164;	// matmul/matmul-hw.mlir:16115:22
  wire [31:0]     a_i_k_8_i_j_3;	// matmul/matmul-hw.mlir:16127:22
  wire [31:0]     b_i_k_8_i_j_3;	// matmul/matmul-hw.mlir:16130:22
  wire [31:0]     c_prev_i_k_8_i_j_3;	// matmul/matmul-hw.mlir:16133:27
  wire            tk_i_k_8_i_j_3;	// matmul/matmul-hw.mlir:16136:23
  wire [31:0]     c_i_k_8_i_j_3;	// matmul/matmul-hw.mlir:16140:22
  reg  [3:0]      i_k_next_3167;	// matmul/matmul-hw.mlir:16145:22
  wire [31:0]     a_i_k_9_i_j_3;	// matmul/matmul-hw.mlir:16157:22
  wire [31:0]     b_i_k_9_i_j_3;	// matmul/matmul-hw.mlir:16160:22
  wire [31:0]     c_prev_i_k_9_i_j_3;	// matmul/matmul-hw.mlir:16163:27
  wire            tk_i_k_9_i_j_3;	// matmul/matmul-hw.mlir:16166:23
  wire [31:0]     c_i_k_9_i_j_3;	// matmul/matmul-hw.mlir:16170:22
  reg  [3:0]      i_k_next_3170;	// matmul/matmul-hw.mlir:16175:22
  wire [31:0]     a_i_k_10_i_j_3;	// matmul/matmul-hw.mlir:16187:23
  wire [31:0]     b_i_k_10_i_j_3;	// matmul/matmul-hw.mlir:16190:23
  wire [31:0]     c_prev_i_k_10_i_j_3;	// matmul/matmul-hw.mlir:16193:28
  wire            tk_i_k_10_i_j_3;	// matmul/matmul-hw.mlir:16196:24
  wire [31:0]     c_i_k_10_i_j_3;	// matmul/matmul-hw.mlir:16200:23
  reg  [3:0]      i_k_next_3173;	// matmul/matmul-hw.mlir:16205:22
  wire [31:0]     a_i_k_11_i_j_3;	// matmul/matmul-hw.mlir:16217:23
  wire [31:0]     b_i_k_11_i_j_3;	// matmul/matmul-hw.mlir:16220:23
  wire [31:0]     c_prev_i_k_11_i_j_3;	// matmul/matmul-hw.mlir:16223:28
  wire            tk_i_k_11_i_j_3;	// matmul/matmul-hw.mlir:16226:24
  wire [31:0]     c_i_k_11_i_j_3;	// matmul/matmul-hw.mlir:16230:23
  reg  [3:0]      i_k_next_3176;	// matmul/matmul-hw.mlir:16235:22
  wire [31:0]     a_i_k_12_i_j_3;	// matmul/matmul-hw.mlir:16247:23
  wire [31:0]     b_i_k_12_i_j_3;	// matmul/matmul-hw.mlir:16250:23
  wire [31:0]     c_prev_i_k_12_i_j_3;	// matmul/matmul-hw.mlir:16253:28
  wire            tk_i_k_12_i_j_3;	// matmul/matmul-hw.mlir:16256:24
  wire [31:0]     c_i_k_12_i_j_3;	// matmul/matmul-hw.mlir:16260:23
  reg  [3:0]      i_k_next_3179;	// matmul/matmul-hw.mlir:16265:22
  wire [31:0]     a_i_k_13_i_j_3;	// matmul/matmul-hw.mlir:16277:23
  wire [31:0]     b_i_k_13_i_j_3;	// matmul/matmul-hw.mlir:16280:23
  wire [31:0]     c_prev_i_k_13_i_j_3;	// matmul/matmul-hw.mlir:16283:28
  wire            tk_i_k_13_i_j_3;	// matmul/matmul-hw.mlir:16286:24
  wire [31:0]     c_i_k_13_i_j_3;	// matmul/matmul-hw.mlir:16290:23
  reg  [3:0]      i_k_next_3182;	// matmul/matmul-hw.mlir:16295:22
  wire [31:0]     a_i_k_14_i_j_3;	// matmul/matmul-hw.mlir:16307:23
  wire [31:0]     b_i_k_14_i_j_3;	// matmul/matmul-hw.mlir:16310:23
  wire [31:0]     c_prev_i_k_14_i_j_3;	// matmul/matmul-hw.mlir:16313:28
  wire            tk_i_k_14_i_j_3;	// matmul/matmul-hw.mlir:16316:24
  wire [31:0]     c_i_k_14_i_j_3;	// matmul/matmul-hw.mlir:16320:23
  reg  [3:0]      i_k_next_3185;	// matmul/matmul-hw.mlir:16325:22
  wire [31:0]     a_i_k_15_i_j_3;	// matmul/matmul-hw.mlir:16337:23
  wire [31:0]     b_i_k_15_i_j_3;	// matmul/matmul-hw.mlir:16340:23
  wire [31:0]     c_prev_i_k_15_i_j_3;	// matmul/matmul-hw.mlir:16343:28
  wire            tk_i_k_15_i_j_3;	// matmul/matmul-hw.mlir:16346:24
  wire [31:0]     c_i_k_15_i_j_3;	// matmul/matmul-hw.mlir:16350:23
  reg  [3:0]      i_k_next_3188;	// matmul/matmul-hw.mlir:16355:22
  reg  [3:0][3:0] i_delayed_3190;	// matmul/matmul-hw.mlir:16364:23
  reg  [3:0]      i_j_next_3194;	// matmul/matmul-hw.mlir:16383:22
  wire [31:0]     a_i_k_0_i_j_4;	// matmul/matmul-hw.mlir:16482:22
  wire [31:0]     b_i_k_0_i_j_4;	// matmul/matmul-hw.mlir:16485:22
  wire [31:0]     c_prev_i_k_0_i_j_4;	// matmul/matmul-hw.mlir:16488:27
  wire            tk_i_k_0_i_j_4;	// matmul/matmul-hw.mlir:16491:23
  wire [31:0]     c_i_k_0_i_j_4;	// matmul/matmul-hw.mlir:16495:22
  reg  [3:0]      i_k_next_3214;	// matmul/matmul-hw.mlir:16500:22
  wire [31:0]     a_i_k_1_i_j_4;	// matmul/matmul-hw.mlir:16512:22
  wire [31:0]     b_i_k_1_i_j_4;	// matmul/matmul-hw.mlir:16515:22
  wire [31:0]     c_prev_i_k_1_i_j_4;	// matmul/matmul-hw.mlir:16518:27
  wire            tk_i_k_1_i_j_4;	// matmul/matmul-hw.mlir:16521:23
  wire [31:0]     c_i_k_1_i_j_4;	// matmul/matmul-hw.mlir:16525:22
  reg  [3:0]      i_k_next_3217;	// matmul/matmul-hw.mlir:16530:22
  wire [31:0]     a_i_k_2_i_j_4;	// matmul/matmul-hw.mlir:16542:22
  wire [31:0]     b_i_k_2_i_j_4;	// matmul/matmul-hw.mlir:16545:22
  wire [31:0]     c_prev_i_k_2_i_j_4;	// matmul/matmul-hw.mlir:16548:27
  wire            tk_i_k_2_i_j_4;	// matmul/matmul-hw.mlir:16551:23
  wire [31:0]     c_i_k_2_i_j_4;	// matmul/matmul-hw.mlir:16555:22
  reg  [3:0]      i_k_next_3220;	// matmul/matmul-hw.mlir:16560:22
  wire [31:0]     a_i_k_3_i_j_4;	// matmul/matmul-hw.mlir:16572:22
  wire [31:0]     b_i_k_3_i_j_4;	// matmul/matmul-hw.mlir:16575:22
  wire [31:0]     c_prev_i_k_3_i_j_4;	// matmul/matmul-hw.mlir:16578:27
  wire            tk_i_k_3_i_j_4;	// matmul/matmul-hw.mlir:16581:23
  wire [31:0]     c_i_k_3_i_j_4;	// matmul/matmul-hw.mlir:16585:22
  reg  [3:0]      i_k_next_3223;	// matmul/matmul-hw.mlir:16590:22
  wire [31:0]     a_i_k_4_i_j_4;	// matmul/matmul-hw.mlir:16602:22
  wire [31:0]     b_i_k_4_i_j_4;	// matmul/matmul-hw.mlir:16605:22
  wire [31:0]     c_prev_i_k_4_i_j_4;	// matmul/matmul-hw.mlir:16608:27
  wire            tk_i_k_4_i_j_4;	// matmul/matmul-hw.mlir:16611:23
  wire [31:0]     c_i_k_4_i_j_4;	// matmul/matmul-hw.mlir:16615:22
  reg  [3:0]      i_k_next_3226;	// matmul/matmul-hw.mlir:16620:22
  wire [31:0]     a_i_k_5_i_j_4;	// matmul/matmul-hw.mlir:16632:22
  wire [31:0]     b_i_k_5_i_j_4;	// matmul/matmul-hw.mlir:16635:22
  wire [31:0]     c_prev_i_k_5_i_j_4;	// matmul/matmul-hw.mlir:16638:27
  wire            tk_i_k_5_i_j_4;	// matmul/matmul-hw.mlir:16641:23
  wire [31:0]     c_i_k_5_i_j_4;	// matmul/matmul-hw.mlir:16645:22
  reg  [3:0]      i_k_next_3229;	// matmul/matmul-hw.mlir:16650:22
  wire [31:0]     a_i_k_6_i_j_4;	// matmul/matmul-hw.mlir:16662:22
  wire [31:0]     b_i_k_6_i_j_4;	// matmul/matmul-hw.mlir:16665:22
  wire [31:0]     c_prev_i_k_6_i_j_4;	// matmul/matmul-hw.mlir:16668:27
  wire            tk_i_k_6_i_j_4;	// matmul/matmul-hw.mlir:16671:23
  wire [31:0]     c_i_k_6_i_j_4;	// matmul/matmul-hw.mlir:16675:22
  reg  [3:0]      i_k_next_3232;	// matmul/matmul-hw.mlir:16680:22
  wire [31:0]     a_i_k_7_i_j_4;	// matmul/matmul-hw.mlir:16692:22
  wire [31:0]     b_i_k_7_i_j_4;	// matmul/matmul-hw.mlir:16695:22
  wire [31:0]     c_prev_i_k_7_i_j_4;	// matmul/matmul-hw.mlir:16698:27
  wire            tk_i_k_7_i_j_4;	// matmul/matmul-hw.mlir:16701:23
  wire [31:0]     c_i_k_7_i_j_4;	// matmul/matmul-hw.mlir:16705:22
  reg  [3:0]      i_k_next_3235;	// matmul/matmul-hw.mlir:16710:22
  wire [31:0]     a_i_k_8_i_j_4;	// matmul/matmul-hw.mlir:16722:22
  wire [31:0]     b_i_k_8_i_j_4;	// matmul/matmul-hw.mlir:16725:22
  wire [31:0]     c_prev_i_k_8_i_j_4;	// matmul/matmul-hw.mlir:16728:27
  wire            tk_i_k_8_i_j_4;	// matmul/matmul-hw.mlir:16731:23
  wire [31:0]     c_i_k_8_i_j_4;	// matmul/matmul-hw.mlir:16735:22
  reg  [3:0]      i_k_next_3238;	// matmul/matmul-hw.mlir:16740:22
  wire [31:0]     a_i_k_9_i_j_4;	// matmul/matmul-hw.mlir:16752:22
  wire [31:0]     b_i_k_9_i_j_4;	// matmul/matmul-hw.mlir:16755:22
  wire [31:0]     c_prev_i_k_9_i_j_4;	// matmul/matmul-hw.mlir:16758:27
  wire            tk_i_k_9_i_j_4;	// matmul/matmul-hw.mlir:16761:23
  wire [31:0]     c_i_k_9_i_j_4;	// matmul/matmul-hw.mlir:16765:22
  reg  [3:0]      i_k_next_3241;	// matmul/matmul-hw.mlir:16770:22
  wire [31:0]     a_i_k_10_i_j_4;	// matmul/matmul-hw.mlir:16782:23
  wire [31:0]     b_i_k_10_i_j_4;	// matmul/matmul-hw.mlir:16785:23
  wire [31:0]     c_prev_i_k_10_i_j_4;	// matmul/matmul-hw.mlir:16788:28
  wire            tk_i_k_10_i_j_4;	// matmul/matmul-hw.mlir:16791:24
  wire [31:0]     c_i_k_10_i_j_4;	// matmul/matmul-hw.mlir:16795:23
  reg  [3:0]      i_k_next_3244;	// matmul/matmul-hw.mlir:16800:22
  wire [31:0]     a_i_k_11_i_j_4;	// matmul/matmul-hw.mlir:16812:23
  wire [31:0]     b_i_k_11_i_j_4;	// matmul/matmul-hw.mlir:16815:23
  wire [31:0]     c_prev_i_k_11_i_j_4;	// matmul/matmul-hw.mlir:16818:28
  wire            tk_i_k_11_i_j_4;	// matmul/matmul-hw.mlir:16821:24
  wire [31:0]     c_i_k_11_i_j_4;	// matmul/matmul-hw.mlir:16825:23
  reg  [3:0]      i_k_next_3247;	// matmul/matmul-hw.mlir:16830:22
  wire [31:0]     a_i_k_12_i_j_4;	// matmul/matmul-hw.mlir:16842:23
  wire [31:0]     b_i_k_12_i_j_4;	// matmul/matmul-hw.mlir:16845:23
  wire [31:0]     c_prev_i_k_12_i_j_4;	// matmul/matmul-hw.mlir:16848:28
  wire            tk_i_k_12_i_j_4;	// matmul/matmul-hw.mlir:16851:24
  wire [31:0]     c_i_k_12_i_j_4;	// matmul/matmul-hw.mlir:16855:23
  reg  [3:0]      i_k_next_3250;	// matmul/matmul-hw.mlir:16860:22
  wire [31:0]     a_i_k_13_i_j_4;	// matmul/matmul-hw.mlir:16872:23
  wire [31:0]     b_i_k_13_i_j_4;	// matmul/matmul-hw.mlir:16875:23
  wire [31:0]     c_prev_i_k_13_i_j_4;	// matmul/matmul-hw.mlir:16878:28
  wire            tk_i_k_13_i_j_4;	// matmul/matmul-hw.mlir:16881:24
  wire [31:0]     c_i_k_13_i_j_4;	// matmul/matmul-hw.mlir:16885:23
  reg  [3:0]      i_k_next_3253;	// matmul/matmul-hw.mlir:16890:22
  wire [31:0]     a_i_k_14_i_j_4;	// matmul/matmul-hw.mlir:16902:23
  wire [31:0]     b_i_k_14_i_j_4;	// matmul/matmul-hw.mlir:16905:23
  wire [31:0]     c_prev_i_k_14_i_j_4;	// matmul/matmul-hw.mlir:16908:28
  wire            tk_i_k_14_i_j_4;	// matmul/matmul-hw.mlir:16911:24
  wire [31:0]     c_i_k_14_i_j_4;	// matmul/matmul-hw.mlir:16915:23
  reg  [3:0]      i_k_next_3256;	// matmul/matmul-hw.mlir:16920:22
  wire [31:0]     a_i_k_15_i_j_4;	// matmul/matmul-hw.mlir:16932:23
  wire [31:0]     b_i_k_15_i_j_4;	// matmul/matmul-hw.mlir:16935:23
  wire [31:0]     c_prev_i_k_15_i_j_4;	// matmul/matmul-hw.mlir:16938:28
  wire            tk_i_k_15_i_j_4;	// matmul/matmul-hw.mlir:16941:24
  wire [31:0]     c_i_k_15_i_j_4;	// matmul/matmul-hw.mlir:16945:23
  reg  [3:0]      i_k_next_3259;	// matmul/matmul-hw.mlir:16950:22
  reg  [3:0][3:0] i_delayed_3261;	// matmul/matmul-hw.mlir:16959:23
  reg  [3:0]      i_j_next_3265;	// matmul/matmul-hw.mlir:16978:22
  wire [31:0]     a_i_k_0_i_j_5;	// matmul/matmul-hw.mlir:17077:22
  wire [31:0]     b_i_k_0_i_j_5;	// matmul/matmul-hw.mlir:17080:22
  wire [31:0]     c_prev_i_k_0_i_j_5;	// matmul/matmul-hw.mlir:17083:27
  wire            tk_i_k_0_i_j_5;	// matmul/matmul-hw.mlir:17086:23
  wire [31:0]     c_i_k_0_i_j_5;	// matmul/matmul-hw.mlir:17090:22
  reg  [3:0]      i_k_next_3285;	// matmul/matmul-hw.mlir:17095:22
  wire [31:0]     a_i_k_1_i_j_5;	// matmul/matmul-hw.mlir:17107:22
  wire [31:0]     b_i_k_1_i_j_5;	// matmul/matmul-hw.mlir:17110:22
  wire [31:0]     c_prev_i_k_1_i_j_5;	// matmul/matmul-hw.mlir:17113:27
  wire            tk_i_k_1_i_j_5;	// matmul/matmul-hw.mlir:17116:23
  wire [31:0]     c_i_k_1_i_j_5;	// matmul/matmul-hw.mlir:17120:22
  reg  [3:0]      i_k_next_3288;	// matmul/matmul-hw.mlir:17125:22
  wire [31:0]     a_i_k_2_i_j_5;	// matmul/matmul-hw.mlir:17137:22
  wire [31:0]     b_i_k_2_i_j_5;	// matmul/matmul-hw.mlir:17140:22
  wire [31:0]     c_prev_i_k_2_i_j_5;	// matmul/matmul-hw.mlir:17143:27
  wire            tk_i_k_2_i_j_5;	// matmul/matmul-hw.mlir:17146:23
  wire [31:0]     c_i_k_2_i_j_5;	// matmul/matmul-hw.mlir:17150:22
  reg  [3:0]      i_k_next_3291;	// matmul/matmul-hw.mlir:17155:22
  wire [31:0]     a_i_k_3_i_j_5;	// matmul/matmul-hw.mlir:17167:22
  wire [31:0]     b_i_k_3_i_j_5;	// matmul/matmul-hw.mlir:17170:22
  wire [31:0]     c_prev_i_k_3_i_j_5;	// matmul/matmul-hw.mlir:17173:27
  wire            tk_i_k_3_i_j_5;	// matmul/matmul-hw.mlir:17176:23
  wire [31:0]     c_i_k_3_i_j_5;	// matmul/matmul-hw.mlir:17180:22
  reg  [3:0]      i_k_next_3294;	// matmul/matmul-hw.mlir:17185:22
  wire [31:0]     a_i_k_4_i_j_5;	// matmul/matmul-hw.mlir:17197:22
  wire [31:0]     b_i_k_4_i_j_5;	// matmul/matmul-hw.mlir:17200:22
  wire [31:0]     c_prev_i_k_4_i_j_5;	// matmul/matmul-hw.mlir:17203:27
  wire            tk_i_k_4_i_j_5;	// matmul/matmul-hw.mlir:17206:23
  wire [31:0]     c_i_k_4_i_j_5;	// matmul/matmul-hw.mlir:17210:22
  reg  [3:0]      i_k_next_3297;	// matmul/matmul-hw.mlir:17215:22
  wire [31:0]     a_i_k_5_i_j_5;	// matmul/matmul-hw.mlir:17227:22
  wire [31:0]     b_i_k_5_i_j_5;	// matmul/matmul-hw.mlir:17230:22
  wire [31:0]     c_prev_i_k_5_i_j_5;	// matmul/matmul-hw.mlir:17233:27
  wire            tk_i_k_5_i_j_5;	// matmul/matmul-hw.mlir:17236:23
  wire [31:0]     c_i_k_5_i_j_5;	// matmul/matmul-hw.mlir:17240:22
  reg  [3:0]      i_k_next_3300;	// matmul/matmul-hw.mlir:17245:22
  wire [31:0]     a_i_k_6_i_j_5;	// matmul/matmul-hw.mlir:17257:22
  wire [31:0]     b_i_k_6_i_j_5;	// matmul/matmul-hw.mlir:17260:22
  wire [31:0]     c_prev_i_k_6_i_j_5;	// matmul/matmul-hw.mlir:17263:27
  wire            tk_i_k_6_i_j_5;	// matmul/matmul-hw.mlir:17266:23
  wire [31:0]     c_i_k_6_i_j_5;	// matmul/matmul-hw.mlir:17270:22
  reg  [3:0]      i_k_next_3303;	// matmul/matmul-hw.mlir:17275:22
  wire [31:0]     a_i_k_7_i_j_5;	// matmul/matmul-hw.mlir:17287:22
  wire [31:0]     b_i_k_7_i_j_5;	// matmul/matmul-hw.mlir:17290:22
  wire [31:0]     c_prev_i_k_7_i_j_5;	// matmul/matmul-hw.mlir:17293:27
  wire            tk_i_k_7_i_j_5;	// matmul/matmul-hw.mlir:17296:23
  wire [31:0]     c_i_k_7_i_j_5;	// matmul/matmul-hw.mlir:17300:22
  reg  [3:0]      i_k_next_3306;	// matmul/matmul-hw.mlir:17305:22
  wire [31:0]     a_i_k_8_i_j_5;	// matmul/matmul-hw.mlir:17317:22
  wire [31:0]     b_i_k_8_i_j_5;	// matmul/matmul-hw.mlir:17320:22
  wire [31:0]     c_prev_i_k_8_i_j_5;	// matmul/matmul-hw.mlir:17323:27
  wire            tk_i_k_8_i_j_5;	// matmul/matmul-hw.mlir:17326:23
  wire [31:0]     c_i_k_8_i_j_5;	// matmul/matmul-hw.mlir:17330:22
  reg  [3:0]      i_k_next_3309;	// matmul/matmul-hw.mlir:17335:22
  wire [31:0]     a_i_k_9_i_j_5;	// matmul/matmul-hw.mlir:17347:22
  wire [31:0]     b_i_k_9_i_j_5;	// matmul/matmul-hw.mlir:17350:22
  wire [31:0]     c_prev_i_k_9_i_j_5;	// matmul/matmul-hw.mlir:17353:27
  wire            tk_i_k_9_i_j_5;	// matmul/matmul-hw.mlir:17356:23
  wire [31:0]     c_i_k_9_i_j_5;	// matmul/matmul-hw.mlir:17360:22
  reg  [3:0]      i_k_next_3312;	// matmul/matmul-hw.mlir:17365:22
  wire [31:0]     a_i_k_10_i_j_5;	// matmul/matmul-hw.mlir:17377:23
  wire [31:0]     b_i_k_10_i_j_5;	// matmul/matmul-hw.mlir:17380:23
  wire [31:0]     c_prev_i_k_10_i_j_5;	// matmul/matmul-hw.mlir:17383:28
  wire            tk_i_k_10_i_j_5;	// matmul/matmul-hw.mlir:17386:24
  wire [31:0]     c_i_k_10_i_j_5;	// matmul/matmul-hw.mlir:17390:23
  reg  [3:0]      i_k_next_3315;	// matmul/matmul-hw.mlir:17395:22
  wire [31:0]     a_i_k_11_i_j_5;	// matmul/matmul-hw.mlir:17407:23
  wire [31:0]     b_i_k_11_i_j_5;	// matmul/matmul-hw.mlir:17410:23
  wire [31:0]     c_prev_i_k_11_i_j_5;	// matmul/matmul-hw.mlir:17413:28
  wire            tk_i_k_11_i_j_5;	// matmul/matmul-hw.mlir:17416:24
  wire [31:0]     c_i_k_11_i_j_5;	// matmul/matmul-hw.mlir:17420:23
  reg  [3:0]      i_k_next_3318;	// matmul/matmul-hw.mlir:17425:22
  wire [31:0]     a_i_k_12_i_j_5;	// matmul/matmul-hw.mlir:17437:23
  wire [31:0]     b_i_k_12_i_j_5;	// matmul/matmul-hw.mlir:17440:23
  wire [31:0]     c_prev_i_k_12_i_j_5;	// matmul/matmul-hw.mlir:17443:28
  wire            tk_i_k_12_i_j_5;	// matmul/matmul-hw.mlir:17446:24
  wire [31:0]     c_i_k_12_i_j_5;	// matmul/matmul-hw.mlir:17450:23
  reg  [3:0]      i_k_next_3321;	// matmul/matmul-hw.mlir:17455:22
  wire [31:0]     a_i_k_13_i_j_5;	// matmul/matmul-hw.mlir:17467:23
  wire [31:0]     b_i_k_13_i_j_5;	// matmul/matmul-hw.mlir:17470:23
  wire [31:0]     c_prev_i_k_13_i_j_5;	// matmul/matmul-hw.mlir:17473:28
  wire            tk_i_k_13_i_j_5;	// matmul/matmul-hw.mlir:17476:24
  wire [31:0]     c_i_k_13_i_j_5;	// matmul/matmul-hw.mlir:17480:23
  reg  [3:0]      i_k_next_3324;	// matmul/matmul-hw.mlir:17485:22
  wire [31:0]     a_i_k_14_i_j_5;	// matmul/matmul-hw.mlir:17497:23
  wire [31:0]     b_i_k_14_i_j_5;	// matmul/matmul-hw.mlir:17500:23
  wire [31:0]     c_prev_i_k_14_i_j_5;	// matmul/matmul-hw.mlir:17503:28
  wire            tk_i_k_14_i_j_5;	// matmul/matmul-hw.mlir:17506:24
  wire [31:0]     c_i_k_14_i_j_5;	// matmul/matmul-hw.mlir:17510:23
  reg  [3:0]      i_k_next_3327;	// matmul/matmul-hw.mlir:17515:22
  wire [31:0]     a_i_k_15_i_j_5;	// matmul/matmul-hw.mlir:17527:23
  wire [31:0]     b_i_k_15_i_j_5;	// matmul/matmul-hw.mlir:17530:23
  wire [31:0]     c_prev_i_k_15_i_j_5;	// matmul/matmul-hw.mlir:17533:28
  wire            tk_i_k_15_i_j_5;	// matmul/matmul-hw.mlir:17536:24
  wire [31:0]     c_i_k_15_i_j_5;	// matmul/matmul-hw.mlir:17540:23
  reg  [3:0]      i_k_next_3330;	// matmul/matmul-hw.mlir:17545:22
  reg  [3:0][3:0] i_delayed_3332;	// matmul/matmul-hw.mlir:17554:23
  reg  [3:0]      i_j_next_3336;	// matmul/matmul-hw.mlir:17573:22
  wire [31:0]     a_i_k_0_i_j_6;	// matmul/matmul-hw.mlir:17672:22
  wire [31:0]     b_i_k_0_i_j_6;	// matmul/matmul-hw.mlir:17675:22
  wire [31:0]     c_prev_i_k_0_i_j_6;	// matmul/matmul-hw.mlir:17678:27
  wire            tk_i_k_0_i_j_6;	// matmul/matmul-hw.mlir:17681:23
  wire [31:0]     c_i_k_0_i_j_6;	// matmul/matmul-hw.mlir:17685:22
  reg  [3:0]      i_k_next_3356;	// matmul/matmul-hw.mlir:17690:22
  wire [31:0]     a_i_k_1_i_j_6;	// matmul/matmul-hw.mlir:17702:22
  wire [31:0]     b_i_k_1_i_j_6;	// matmul/matmul-hw.mlir:17705:22
  wire [31:0]     c_prev_i_k_1_i_j_6;	// matmul/matmul-hw.mlir:17708:27
  wire            tk_i_k_1_i_j_6;	// matmul/matmul-hw.mlir:17711:23
  wire [31:0]     c_i_k_1_i_j_6;	// matmul/matmul-hw.mlir:17715:22
  reg  [3:0]      i_k_next_3359;	// matmul/matmul-hw.mlir:17720:22
  wire [31:0]     a_i_k_2_i_j_6;	// matmul/matmul-hw.mlir:17732:22
  wire [31:0]     b_i_k_2_i_j_6;	// matmul/matmul-hw.mlir:17735:22
  wire [31:0]     c_prev_i_k_2_i_j_6;	// matmul/matmul-hw.mlir:17738:27
  wire            tk_i_k_2_i_j_6;	// matmul/matmul-hw.mlir:17741:23
  wire [31:0]     c_i_k_2_i_j_6;	// matmul/matmul-hw.mlir:17745:22
  reg  [3:0]      i_k_next_3362;	// matmul/matmul-hw.mlir:17750:22
  wire [31:0]     a_i_k_3_i_j_6;	// matmul/matmul-hw.mlir:17762:22
  wire [31:0]     b_i_k_3_i_j_6;	// matmul/matmul-hw.mlir:17765:22
  wire [31:0]     c_prev_i_k_3_i_j_6;	// matmul/matmul-hw.mlir:17768:27
  wire            tk_i_k_3_i_j_6;	// matmul/matmul-hw.mlir:17771:23
  wire [31:0]     c_i_k_3_i_j_6;	// matmul/matmul-hw.mlir:17775:22
  reg  [3:0]      i_k_next_3365;	// matmul/matmul-hw.mlir:17780:22
  wire [31:0]     a_i_k_4_i_j_6;	// matmul/matmul-hw.mlir:17792:22
  wire [31:0]     b_i_k_4_i_j_6;	// matmul/matmul-hw.mlir:17795:22
  wire [31:0]     c_prev_i_k_4_i_j_6;	// matmul/matmul-hw.mlir:17798:27
  wire            tk_i_k_4_i_j_6;	// matmul/matmul-hw.mlir:17801:23
  wire [31:0]     c_i_k_4_i_j_6;	// matmul/matmul-hw.mlir:17805:22
  reg  [3:0]      i_k_next_3368;	// matmul/matmul-hw.mlir:17810:22
  wire [31:0]     a_i_k_5_i_j_6;	// matmul/matmul-hw.mlir:17822:22
  wire [31:0]     b_i_k_5_i_j_6;	// matmul/matmul-hw.mlir:17825:22
  wire [31:0]     c_prev_i_k_5_i_j_6;	// matmul/matmul-hw.mlir:17828:27
  wire            tk_i_k_5_i_j_6;	// matmul/matmul-hw.mlir:17831:23
  wire [31:0]     c_i_k_5_i_j_6;	// matmul/matmul-hw.mlir:17835:22
  reg  [3:0]      i_k_next_3371;	// matmul/matmul-hw.mlir:17840:22
  wire [31:0]     a_i_k_6_i_j_6;	// matmul/matmul-hw.mlir:17852:22
  wire [31:0]     b_i_k_6_i_j_6;	// matmul/matmul-hw.mlir:17855:22
  wire [31:0]     c_prev_i_k_6_i_j_6;	// matmul/matmul-hw.mlir:17858:27
  wire            tk_i_k_6_i_j_6;	// matmul/matmul-hw.mlir:17861:23
  wire [31:0]     c_i_k_6_i_j_6;	// matmul/matmul-hw.mlir:17865:22
  reg  [3:0]      i_k_next_3374;	// matmul/matmul-hw.mlir:17870:22
  wire [31:0]     a_i_k_7_i_j_6;	// matmul/matmul-hw.mlir:17882:22
  wire [31:0]     b_i_k_7_i_j_6;	// matmul/matmul-hw.mlir:17885:22
  wire [31:0]     c_prev_i_k_7_i_j_6;	// matmul/matmul-hw.mlir:17888:27
  wire            tk_i_k_7_i_j_6;	// matmul/matmul-hw.mlir:17891:23
  wire [31:0]     c_i_k_7_i_j_6;	// matmul/matmul-hw.mlir:17895:22
  reg  [3:0]      i_k_next_3377;	// matmul/matmul-hw.mlir:17900:22
  wire [31:0]     a_i_k_8_i_j_6;	// matmul/matmul-hw.mlir:17912:22
  wire [31:0]     b_i_k_8_i_j_6;	// matmul/matmul-hw.mlir:17915:22
  wire [31:0]     c_prev_i_k_8_i_j_6;	// matmul/matmul-hw.mlir:17918:27
  wire            tk_i_k_8_i_j_6;	// matmul/matmul-hw.mlir:17921:23
  wire [31:0]     c_i_k_8_i_j_6;	// matmul/matmul-hw.mlir:17925:22
  reg  [3:0]      i_k_next_3380;	// matmul/matmul-hw.mlir:17930:22
  wire [31:0]     a_i_k_9_i_j_6;	// matmul/matmul-hw.mlir:17942:22
  wire [31:0]     b_i_k_9_i_j_6;	// matmul/matmul-hw.mlir:17945:22
  wire [31:0]     c_prev_i_k_9_i_j_6;	// matmul/matmul-hw.mlir:17948:27
  wire            tk_i_k_9_i_j_6;	// matmul/matmul-hw.mlir:17951:23
  wire [31:0]     c_i_k_9_i_j_6;	// matmul/matmul-hw.mlir:17955:22
  reg  [3:0]      i_k_next_3383;	// matmul/matmul-hw.mlir:17960:22
  wire [31:0]     a_i_k_10_i_j_6;	// matmul/matmul-hw.mlir:17972:23
  wire [31:0]     b_i_k_10_i_j_6;	// matmul/matmul-hw.mlir:17975:23
  wire [31:0]     c_prev_i_k_10_i_j_6;	// matmul/matmul-hw.mlir:17978:28
  wire            tk_i_k_10_i_j_6;	// matmul/matmul-hw.mlir:17981:24
  wire [31:0]     c_i_k_10_i_j_6;	// matmul/matmul-hw.mlir:17985:23
  reg  [3:0]      i_k_next_3386;	// matmul/matmul-hw.mlir:17990:22
  wire [31:0]     a_i_k_11_i_j_6;	// matmul/matmul-hw.mlir:18002:23
  wire [31:0]     b_i_k_11_i_j_6;	// matmul/matmul-hw.mlir:18005:23
  wire [31:0]     c_prev_i_k_11_i_j_6;	// matmul/matmul-hw.mlir:18008:28
  wire            tk_i_k_11_i_j_6;	// matmul/matmul-hw.mlir:18011:24
  wire [31:0]     c_i_k_11_i_j_6;	// matmul/matmul-hw.mlir:18015:23
  reg  [3:0]      i_k_next_3389;	// matmul/matmul-hw.mlir:18020:22
  wire [31:0]     a_i_k_12_i_j_6;	// matmul/matmul-hw.mlir:18032:23
  wire [31:0]     b_i_k_12_i_j_6;	// matmul/matmul-hw.mlir:18035:23
  wire [31:0]     c_prev_i_k_12_i_j_6;	// matmul/matmul-hw.mlir:18038:28
  wire            tk_i_k_12_i_j_6;	// matmul/matmul-hw.mlir:18041:24
  wire [31:0]     c_i_k_12_i_j_6;	// matmul/matmul-hw.mlir:18045:23
  reg  [3:0]      i_k_next_3392;	// matmul/matmul-hw.mlir:18050:22
  wire [31:0]     a_i_k_13_i_j_6;	// matmul/matmul-hw.mlir:18062:23
  wire [31:0]     b_i_k_13_i_j_6;	// matmul/matmul-hw.mlir:18065:23
  wire [31:0]     c_prev_i_k_13_i_j_6;	// matmul/matmul-hw.mlir:18068:28
  wire            tk_i_k_13_i_j_6;	// matmul/matmul-hw.mlir:18071:24
  wire [31:0]     c_i_k_13_i_j_6;	// matmul/matmul-hw.mlir:18075:23
  reg  [3:0]      i_k_next_3395;	// matmul/matmul-hw.mlir:18080:22
  wire [31:0]     a_i_k_14_i_j_6;	// matmul/matmul-hw.mlir:18092:23
  wire [31:0]     b_i_k_14_i_j_6;	// matmul/matmul-hw.mlir:18095:23
  wire [31:0]     c_prev_i_k_14_i_j_6;	// matmul/matmul-hw.mlir:18098:28
  wire            tk_i_k_14_i_j_6;	// matmul/matmul-hw.mlir:18101:24
  wire [31:0]     c_i_k_14_i_j_6;	// matmul/matmul-hw.mlir:18105:23
  reg  [3:0]      i_k_next_3398;	// matmul/matmul-hw.mlir:18110:22
  wire [31:0]     a_i_k_15_i_j_6;	// matmul/matmul-hw.mlir:18122:23
  wire [31:0]     b_i_k_15_i_j_6;	// matmul/matmul-hw.mlir:18125:23
  wire [31:0]     c_prev_i_k_15_i_j_6;	// matmul/matmul-hw.mlir:18128:28
  wire            tk_i_k_15_i_j_6;	// matmul/matmul-hw.mlir:18131:24
  wire [31:0]     c_i_k_15_i_j_6;	// matmul/matmul-hw.mlir:18135:23
  reg  [3:0]      i_k_next_3401;	// matmul/matmul-hw.mlir:18140:22
  reg  [3:0][3:0] i_delayed_3403;	// matmul/matmul-hw.mlir:18149:23
  reg  [3:0]      i_j_next_3407;	// matmul/matmul-hw.mlir:18168:22
  wire [31:0]     a_i_k_0_i_j_7;	// matmul/matmul-hw.mlir:18267:22
  wire [31:0]     b_i_k_0_i_j_7;	// matmul/matmul-hw.mlir:18270:22
  wire [31:0]     c_prev_i_k_0_i_j_7;	// matmul/matmul-hw.mlir:18273:27
  wire            tk_i_k_0_i_j_7;	// matmul/matmul-hw.mlir:18276:23
  wire [31:0]     c_i_k_0_i_j_7;	// matmul/matmul-hw.mlir:18280:22
  reg  [3:0]      i_k_next_3427;	// matmul/matmul-hw.mlir:18285:22
  wire [31:0]     a_i_k_1_i_j_7;	// matmul/matmul-hw.mlir:18297:22
  wire [31:0]     b_i_k_1_i_j_7;	// matmul/matmul-hw.mlir:18300:22
  wire [31:0]     c_prev_i_k_1_i_j_7;	// matmul/matmul-hw.mlir:18303:27
  wire            tk_i_k_1_i_j_7;	// matmul/matmul-hw.mlir:18306:23
  wire [31:0]     c_i_k_1_i_j_7;	// matmul/matmul-hw.mlir:18310:22
  reg  [3:0]      i_k_next_3430;	// matmul/matmul-hw.mlir:18315:22
  wire [31:0]     a_i_k_2_i_j_7;	// matmul/matmul-hw.mlir:18327:22
  wire [31:0]     b_i_k_2_i_j_7;	// matmul/matmul-hw.mlir:18330:22
  wire [31:0]     c_prev_i_k_2_i_j_7;	// matmul/matmul-hw.mlir:18333:27
  wire            tk_i_k_2_i_j_7;	// matmul/matmul-hw.mlir:18336:23
  wire [31:0]     c_i_k_2_i_j_7;	// matmul/matmul-hw.mlir:18340:22
  reg  [3:0]      i_k_next_3433;	// matmul/matmul-hw.mlir:18345:22
  wire [31:0]     a_i_k_3_i_j_7;	// matmul/matmul-hw.mlir:18357:22
  wire [31:0]     b_i_k_3_i_j_7;	// matmul/matmul-hw.mlir:18360:22
  wire [31:0]     c_prev_i_k_3_i_j_7;	// matmul/matmul-hw.mlir:18363:27
  wire            tk_i_k_3_i_j_7;	// matmul/matmul-hw.mlir:18366:23
  wire [31:0]     c_i_k_3_i_j_7;	// matmul/matmul-hw.mlir:18370:22
  reg  [3:0]      i_k_next_3436;	// matmul/matmul-hw.mlir:18375:22
  wire [31:0]     a_i_k_4_i_j_7;	// matmul/matmul-hw.mlir:18387:22
  wire [31:0]     b_i_k_4_i_j_7;	// matmul/matmul-hw.mlir:18390:22
  wire [31:0]     c_prev_i_k_4_i_j_7;	// matmul/matmul-hw.mlir:18393:27
  wire            tk_i_k_4_i_j_7;	// matmul/matmul-hw.mlir:18396:23
  wire [31:0]     c_i_k_4_i_j_7;	// matmul/matmul-hw.mlir:18400:22
  reg  [3:0]      i_k_next_3439;	// matmul/matmul-hw.mlir:18405:22
  wire [31:0]     a_i_k_5_i_j_7;	// matmul/matmul-hw.mlir:18417:22
  wire [31:0]     b_i_k_5_i_j_7;	// matmul/matmul-hw.mlir:18420:22
  wire [31:0]     c_prev_i_k_5_i_j_7;	// matmul/matmul-hw.mlir:18423:27
  wire            tk_i_k_5_i_j_7;	// matmul/matmul-hw.mlir:18426:23
  wire [31:0]     c_i_k_5_i_j_7;	// matmul/matmul-hw.mlir:18430:22
  reg  [3:0]      i_k_next_3442;	// matmul/matmul-hw.mlir:18435:22
  wire [31:0]     a_i_k_6_i_j_7;	// matmul/matmul-hw.mlir:18447:22
  wire [31:0]     b_i_k_6_i_j_7;	// matmul/matmul-hw.mlir:18450:22
  wire [31:0]     c_prev_i_k_6_i_j_7;	// matmul/matmul-hw.mlir:18453:27
  wire            tk_i_k_6_i_j_7;	// matmul/matmul-hw.mlir:18456:23
  wire [31:0]     c_i_k_6_i_j_7;	// matmul/matmul-hw.mlir:18460:22
  reg  [3:0]      i_k_next_3445;	// matmul/matmul-hw.mlir:18465:22
  wire [31:0]     a_i_k_7_i_j_7;	// matmul/matmul-hw.mlir:18477:22
  wire [31:0]     b_i_k_7_i_j_7;	// matmul/matmul-hw.mlir:18480:22
  wire [31:0]     c_prev_i_k_7_i_j_7;	// matmul/matmul-hw.mlir:18483:27
  wire            tk_i_k_7_i_j_7;	// matmul/matmul-hw.mlir:18486:23
  wire [31:0]     c_i_k_7_i_j_7;	// matmul/matmul-hw.mlir:18490:22
  reg  [3:0]      i_k_next_3448;	// matmul/matmul-hw.mlir:18495:22
  wire [31:0]     a_i_k_8_i_j_7;	// matmul/matmul-hw.mlir:18507:22
  wire [31:0]     b_i_k_8_i_j_7;	// matmul/matmul-hw.mlir:18510:22
  wire [31:0]     c_prev_i_k_8_i_j_7;	// matmul/matmul-hw.mlir:18513:27
  wire            tk_i_k_8_i_j_7;	// matmul/matmul-hw.mlir:18516:23
  wire [31:0]     c_i_k_8_i_j_7;	// matmul/matmul-hw.mlir:18520:22
  reg  [3:0]      i_k_next_3451;	// matmul/matmul-hw.mlir:18525:22
  wire [31:0]     a_i_k_9_i_j_7;	// matmul/matmul-hw.mlir:18537:22
  wire [31:0]     b_i_k_9_i_j_7;	// matmul/matmul-hw.mlir:18540:22
  wire [31:0]     c_prev_i_k_9_i_j_7;	// matmul/matmul-hw.mlir:18543:27
  wire            tk_i_k_9_i_j_7;	// matmul/matmul-hw.mlir:18546:23
  wire [31:0]     c_i_k_9_i_j_7;	// matmul/matmul-hw.mlir:18550:22
  reg  [3:0]      i_k_next_3454;	// matmul/matmul-hw.mlir:18555:22
  wire [31:0]     a_i_k_10_i_j_7;	// matmul/matmul-hw.mlir:18567:23
  wire [31:0]     b_i_k_10_i_j_7;	// matmul/matmul-hw.mlir:18570:23
  wire [31:0]     c_prev_i_k_10_i_j_7;	// matmul/matmul-hw.mlir:18573:28
  wire            tk_i_k_10_i_j_7;	// matmul/matmul-hw.mlir:18576:24
  wire [31:0]     c_i_k_10_i_j_7;	// matmul/matmul-hw.mlir:18580:23
  reg  [3:0]      i_k_next_3457;	// matmul/matmul-hw.mlir:18585:22
  wire [31:0]     a_i_k_11_i_j_7;	// matmul/matmul-hw.mlir:18597:23
  wire [31:0]     b_i_k_11_i_j_7;	// matmul/matmul-hw.mlir:18600:23
  wire [31:0]     c_prev_i_k_11_i_j_7;	// matmul/matmul-hw.mlir:18603:28
  wire            tk_i_k_11_i_j_7;	// matmul/matmul-hw.mlir:18606:24
  wire [31:0]     c_i_k_11_i_j_7;	// matmul/matmul-hw.mlir:18610:23
  reg  [3:0]      i_k_next_3460;	// matmul/matmul-hw.mlir:18615:22
  wire [31:0]     a_i_k_12_i_j_7;	// matmul/matmul-hw.mlir:18627:23
  wire [31:0]     b_i_k_12_i_j_7;	// matmul/matmul-hw.mlir:18630:23
  wire [31:0]     c_prev_i_k_12_i_j_7;	// matmul/matmul-hw.mlir:18633:28
  wire            tk_i_k_12_i_j_7;	// matmul/matmul-hw.mlir:18636:24
  wire [31:0]     c_i_k_12_i_j_7;	// matmul/matmul-hw.mlir:18640:23
  reg  [3:0]      i_k_next_3463;	// matmul/matmul-hw.mlir:18645:22
  wire [31:0]     a_i_k_13_i_j_7;	// matmul/matmul-hw.mlir:18657:23
  wire [31:0]     b_i_k_13_i_j_7;	// matmul/matmul-hw.mlir:18660:23
  wire [31:0]     c_prev_i_k_13_i_j_7;	// matmul/matmul-hw.mlir:18663:28
  wire            tk_i_k_13_i_j_7;	// matmul/matmul-hw.mlir:18666:24
  wire [31:0]     c_i_k_13_i_j_7;	// matmul/matmul-hw.mlir:18670:23
  reg  [3:0]      i_k_next_3466;	// matmul/matmul-hw.mlir:18675:22
  wire [31:0]     a_i_k_14_i_j_7;	// matmul/matmul-hw.mlir:18687:23
  wire [31:0]     b_i_k_14_i_j_7;	// matmul/matmul-hw.mlir:18690:23
  wire [31:0]     c_prev_i_k_14_i_j_7;	// matmul/matmul-hw.mlir:18693:28
  wire            tk_i_k_14_i_j_7;	// matmul/matmul-hw.mlir:18696:24
  wire [31:0]     c_i_k_14_i_j_7;	// matmul/matmul-hw.mlir:18700:23
  reg  [3:0]      i_k_next_3469;	// matmul/matmul-hw.mlir:18705:22
  wire [31:0]     a_i_k_15_i_j_7;	// matmul/matmul-hw.mlir:18717:23
  wire [31:0]     b_i_k_15_i_j_7;	// matmul/matmul-hw.mlir:18720:23
  wire [31:0]     c_prev_i_k_15_i_j_7;	// matmul/matmul-hw.mlir:18723:28
  wire            tk_i_k_15_i_j_7;	// matmul/matmul-hw.mlir:18726:24
  wire [31:0]     c_i_k_15_i_j_7;	// matmul/matmul-hw.mlir:18730:23
  reg  [3:0]      i_k_next_3472;	// matmul/matmul-hw.mlir:18735:22
  reg  [3:0][3:0] i_delayed_3474;	// matmul/matmul-hw.mlir:18744:23
  reg  [3:0]      i_j_next_3478;	// matmul/matmul-hw.mlir:18763:22
  wire [31:0]     a_i_k_0_i_j_8;	// matmul/matmul-hw.mlir:18862:22
  wire [31:0]     b_i_k_0_i_j_8;	// matmul/matmul-hw.mlir:18865:22
  wire [31:0]     c_prev_i_k_0_i_j_8;	// matmul/matmul-hw.mlir:18868:27
  wire            tk_i_k_0_i_j_8;	// matmul/matmul-hw.mlir:18871:23
  wire [31:0]     c_i_k_0_i_j_8;	// matmul/matmul-hw.mlir:18875:22
  reg  [3:0]      i_k_next_3498;	// matmul/matmul-hw.mlir:18880:22
  wire [31:0]     a_i_k_1_i_j_8;	// matmul/matmul-hw.mlir:18892:22
  wire [31:0]     b_i_k_1_i_j_8;	// matmul/matmul-hw.mlir:18895:22
  wire [31:0]     c_prev_i_k_1_i_j_8;	// matmul/matmul-hw.mlir:18898:27
  wire            tk_i_k_1_i_j_8;	// matmul/matmul-hw.mlir:18901:23
  wire [31:0]     c_i_k_1_i_j_8;	// matmul/matmul-hw.mlir:18905:22
  reg  [3:0]      i_k_next_3501;	// matmul/matmul-hw.mlir:18910:22
  wire [31:0]     a_i_k_2_i_j_8;	// matmul/matmul-hw.mlir:18922:22
  wire [31:0]     b_i_k_2_i_j_8;	// matmul/matmul-hw.mlir:18925:22
  wire [31:0]     c_prev_i_k_2_i_j_8;	// matmul/matmul-hw.mlir:18928:27
  wire            tk_i_k_2_i_j_8;	// matmul/matmul-hw.mlir:18931:23
  wire [31:0]     c_i_k_2_i_j_8;	// matmul/matmul-hw.mlir:18935:22
  reg  [3:0]      i_k_next_3504;	// matmul/matmul-hw.mlir:18940:22
  wire [31:0]     a_i_k_3_i_j_8;	// matmul/matmul-hw.mlir:18952:22
  wire [31:0]     b_i_k_3_i_j_8;	// matmul/matmul-hw.mlir:18955:22
  wire [31:0]     c_prev_i_k_3_i_j_8;	// matmul/matmul-hw.mlir:18958:27
  wire            tk_i_k_3_i_j_8;	// matmul/matmul-hw.mlir:18961:23
  wire [31:0]     c_i_k_3_i_j_8;	// matmul/matmul-hw.mlir:18965:22
  reg  [3:0]      i_k_next_3507;	// matmul/matmul-hw.mlir:18970:22
  wire [31:0]     a_i_k_4_i_j_8;	// matmul/matmul-hw.mlir:18982:22
  wire [31:0]     b_i_k_4_i_j_8;	// matmul/matmul-hw.mlir:18985:22
  wire [31:0]     c_prev_i_k_4_i_j_8;	// matmul/matmul-hw.mlir:18988:27
  wire            tk_i_k_4_i_j_8;	// matmul/matmul-hw.mlir:18991:23
  wire [31:0]     c_i_k_4_i_j_8;	// matmul/matmul-hw.mlir:18995:22
  reg  [3:0]      i_k_next_3510;	// matmul/matmul-hw.mlir:19000:22
  wire [31:0]     a_i_k_5_i_j_8;	// matmul/matmul-hw.mlir:19012:22
  wire [31:0]     b_i_k_5_i_j_8;	// matmul/matmul-hw.mlir:19015:22
  wire [31:0]     c_prev_i_k_5_i_j_8;	// matmul/matmul-hw.mlir:19018:27
  wire            tk_i_k_5_i_j_8;	// matmul/matmul-hw.mlir:19021:23
  wire [31:0]     c_i_k_5_i_j_8;	// matmul/matmul-hw.mlir:19025:22
  reg  [3:0]      i_k_next_3513;	// matmul/matmul-hw.mlir:19030:22
  wire [31:0]     a_i_k_6_i_j_8;	// matmul/matmul-hw.mlir:19042:22
  wire [31:0]     b_i_k_6_i_j_8;	// matmul/matmul-hw.mlir:19045:22
  wire [31:0]     c_prev_i_k_6_i_j_8;	// matmul/matmul-hw.mlir:19048:27
  wire            tk_i_k_6_i_j_8;	// matmul/matmul-hw.mlir:19051:23
  wire [31:0]     c_i_k_6_i_j_8;	// matmul/matmul-hw.mlir:19055:22
  reg  [3:0]      i_k_next_3516;	// matmul/matmul-hw.mlir:19060:22
  wire [31:0]     a_i_k_7_i_j_8;	// matmul/matmul-hw.mlir:19072:22
  wire [31:0]     b_i_k_7_i_j_8;	// matmul/matmul-hw.mlir:19075:22
  wire [31:0]     c_prev_i_k_7_i_j_8;	// matmul/matmul-hw.mlir:19078:27
  wire            tk_i_k_7_i_j_8;	// matmul/matmul-hw.mlir:19081:23
  wire [31:0]     c_i_k_7_i_j_8;	// matmul/matmul-hw.mlir:19085:22
  reg  [3:0]      i_k_next_3519;	// matmul/matmul-hw.mlir:19090:22
  wire [31:0]     a_i_k_8_i_j_8;	// matmul/matmul-hw.mlir:19102:22
  wire [31:0]     b_i_k_8_i_j_8;	// matmul/matmul-hw.mlir:19105:22
  wire [31:0]     c_prev_i_k_8_i_j_8;	// matmul/matmul-hw.mlir:19108:27
  wire            tk_i_k_8_i_j_8;	// matmul/matmul-hw.mlir:19111:23
  wire [31:0]     c_i_k_8_i_j_8;	// matmul/matmul-hw.mlir:19115:22
  reg  [3:0]      i_k_next_3522;	// matmul/matmul-hw.mlir:19120:22
  wire [31:0]     a_i_k_9_i_j_8;	// matmul/matmul-hw.mlir:19132:22
  wire [31:0]     b_i_k_9_i_j_8;	// matmul/matmul-hw.mlir:19135:22
  wire [31:0]     c_prev_i_k_9_i_j_8;	// matmul/matmul-hw.mlir:19138:27
  wire            tk_i_k_9_i_j_8;	// matmul/matmul-hw.mlir:19141:23
  wire [31:0]     c_i_k_9_i_j_8;	// matmul/matmul-hw.mlir:19145:22
  reg  [3:0]      i_k_next_3525;	// matmul/matmul-hw.mlir:19150:22
  wire [31:0]     a_i_k_10_i_j_8;	// matmul/matmul-hw.mlir:19162:23
  wire [31:0]     b_i_k_10_i_j_8;	// matmul/matmul-hw.mlir:19165:23
  wire [31:0]     c_prev_i_k_10_i_j_8;	// matmul/matmul-hw.mlir:19168:28
  wire            tk_i_k_10_i_j_8;	// matmul/matmul-hw.mlir:19171:24
  wire [31:0]     c_i_k_10_i_j_8;	// matmul/matmul-hw.mlir:19175:23
  reg  [3:0]      i_k_next_3528;	// matmul/matmul-hw.mlir:19180:22
  wire [31:0]     a_i_k_11_i_j_8;	// matmul/matmul-hw.mlir:19192:23
  wire [31:0]     b_i_k_11_i_j_8;	// matmul/matmul-hw.mlir:19195:23
  wire [31:0]     c_prev_i_k_11_i_j_8;	// matmul/matmul-hw.mlir:19198:28
  wire            tk_i_k_11_i_j_8;	// matmul/matmul-hw.mlir:19201:24
  wire [31:0]     c_i_k_11_i_j_8;	// matmul/matmul-hw.mlir:19205:23
  reg  [3:0]      i_k_next_3531;	// matmul/matmul-hw.mlir:19210:22
  wire [31:0]     a_i_k_12_i_j_8;	// matmul/matmul-hw.mlir:19222:23
  wire [31:0]     b_i_k_12_i_j_8;	// matmul/matmul-hw.mlir:19225:23
  wire [31:0]     c_prev_i_k_12_i_j_8;	// matmul/matmul-hw.mlir:19228:28
  wire            tk_i_k_12_i_j_8;	// matmul/matmul-hw.mlir:19231:24
  wire [31:0]     c_i_k_12_i_j_8;	// matmul/matmul-hw.mlir:19235:23
  reg  [3:0]      i_k_next_3534;	// matmul/matmul-hw.mlir:19240:22
  wire [31:0]     a_i_k_13_i_j_8;	// matmul/matmul-hw.mlir:19252:23
  wire [31:0]     b_i_k_13_i_j_8;	// matmul/matmul-hw.mlir:19255:23
  wire [31:0]     c_prev_i_k_13_i_j_8;	// matmul/matmul-hw.mlir:19258:28
  wire            tk_i_k_13_i_j_8;	// matmul/matmul-hw.mlir:19261:24
  wire [31:0]     c_i_k_13_i_j_8;	// matmul/matmul-hw.mlir:19265:23
  reg  [3:0]      i_k_next_3537;	// matmul/matmul-hw.mlir:19270:22
  wire [31:0]     a_i_k_14_i_j_8;	// matmul/matmul-hw.mlir:19282:23
  wire [31:0]     b_i_k_14_i_j_8;	// matmul/matmul-hw.mlir:19285:23
  wire [31:0]     c_prev_i_k_14_i_j_8;	// matmul/matmul-hw.mlir:19288:28
  wire            tk_i_k_14_i_j_8;	// matmul/matmul-hw.mlir:19291:24
  wire [31:0]     c_i_k_14_i_j_8;	// matmul/matmul-hw.mlir:19295:23
  reg  [3:0]      i_k_next_3540;	// matmul/matmul-hw.mlir:19300:22
  wire [31:0]     a_i_k_15_i_j_8;	// matmul/matmul-hw.mlir:19312:23
  wire [31:0]     b_i_k_15_i_j_8;	// matmul/matmul-hw.mlir:19315:23
  wire [31:0]     c_prev_i_k_15_i_j_8;	// matmul/matmul-hw.mlir:19318:28
  wire            tk_i_k_15_i_j_8;	// matmul/matmul-hw.mlir:19321:24
  wire [31:0]     c_i_k_15_i_j_8;	// matmul/matmul-hw.mlir:19325:23
  reg  [3:0]      i_k_next_3543;	// matmul/matmul-hw.mlir:19330:22
  reg  [3:0][3:0] i_delayed_3545;	// matmul/matmul-hw.mlir:19339:23
  reg  [3:0]      i_j_next_3549;	// matmul/matmul-hw.mlir:19358:22
  wire [31:0]     a_i_k_0_i_j_9;	// matmul/matmul-hw.mlir:19457:22
  wire [31:0]     b_i_k_0_i_j_9;	// matmul/matmul-hw.mlir:19460:22
  wire [31:0]     c_prev_i_k_0_i_j_9;	// matmul/matmul-hw.mlir:19463:27
  wire            tk_i_k_0_i_j_9;	// matmul/matmul-hw.mlir:19466:23
  wire [31:0]     c_i_k_0_i_j_9;	// matmul/matmul-hw.mlir:19470:22
  reg  [3:0]      i_k_next_3569;	// matmul/matmul-hw.mlir:19475:22
  wire [31:0]     a_i_k_1_i_j_9;	// matmul/matmul-hw.mlir:19487:22
  wire [31:0]     b_i_k_1_i_j_9;	// matmul/matmul-hw.mlir:19490:22
  wire [31:0]     c_prev_i_k_1_i_j_9;	// matmul/matmul-hw.mlir:19493:27
  wire            tk_i_k_1_i_j_9;	// matmul/matmul-hw.mlir:19496:23
  wire [31:0]     c_i_k_1_i_j_9;	// matmul/matmul-hw.mlir:19500:22
  reg  [3:0]      i_k_next_3572;	// matmul/matmul-hw.mlir:19505:22
  wire [31:0]     a_i_k_2_i_j_9;	// matmul/matmul-hw.mlir:19517:22
  wire [31:0]     b_i_k_2_i_j_9;	// matmul/matmul-hw.mlir:19520:22
  wire [31:0]     c_prev_i_k_2_i_j_9;	// matmul/matmul-hw.mlir:19523:27
  wire            tk_i_k_2_i_j_9;	// matmul/matmul-hw.mlir:19526:23
  wire [31:0]     c_i_k_2_i_j_9;	// matmul/matmul-hw.mlir:19530:22
  reg  [3:0]      i_k_next_3575;	// matmul/matmul-hw.mlir:19535:22
  wire [31:0]     a_i_k_3_i_j_9;	// matmul/matmul-hw.mlir:19547:22
  wire [31:0]     b_i_k_3_i_j_9;	// matmul/matmul-hw.mlir:19550:22
  wire [31:0]     c_prev_i_k_3_i_j_9;	// matmul/matmul-hw.mlir:19553:27
  wire            tk_i_k_3_i_j_9;	// matmul/matmul-hw.mlir:19556:23
  wire [31:0]     c_i_k_3_i_j_9;	// matmul/matmul-hw.mlir:19560:22
  reg  [3:0]      i_k_next_3578;	// matmul/matmul-hw.mlir:19565:22
  wire [31:0]     a_i_k_4_i_j_9;	// matmul/matmul-hw.mlir:19577:22
  wire [31:0]     b_i_k_4_i_j_9;	// matmul/matmul-hw.mlir:19580:22
  wire [31:0]     c_prev_i_k_4_i_j_9;	// matmul/matmul-hw.mlir:19583:27
  wire            tk_i_k_4_i_j_9;	// matmul/matmul-hw.mlir:19586:23
  wire [31:0]     c_i_k_4_i_j_9;	// matmul/matmul-hw.mlir:19590:22
  reg  [3:0]      i_k_next_3581;	// matmul/matmul-hw.mlir:19595:22
  wire [31:0]     a_i_k_5_i_j_9;	// matmul/matmul-hw.mlir:19607:22
  wire [31:0]     b_i_k_5_i_j_9;	// matmul/matmul-hw.mlir:19610:22
  wire [31:0]     c_prev_i_k_5_i_j_9;	// matmul/matmul-hw.mlir:19613:27
  wire            tk_i_k_5_i_j_9;	// matmul/matmul-hw.mlir:19616:23
  wire [31:0]     c_i_k_5_i_j_9;	// matmul/matmul-hw.mlir:19620:22
  reg  [3:0]      i_k_next_3584;	// matmul/matmul-hw.mlir:19625:22
  wire [31:0]     a_i_k_6_i_j_9;	// matmul/matmul-hw.mlir:19637:22
  wire [31:0]     b_i_k_6_i_j_9;	// matmul/matmul-hw.mlir:19640:22
  wire [31:0]     c_prev_i_k_6_i_j_9;	// matmul/matmul-hw.mlir:19643:27
  wire            tk_i_k_6_i_j_9;	// matmul/matmul-hw.mlir:19646:23
  wire [31:0]     c_i_k_6_i_j_9;	// matmul/matmul-hw.mlir:19650:22
  reg  [3:0]      i_k_next_3587;	// matmul/matmul-hw.mlir:19655:22
  wire [31:0]     a_i_k_7_i_j_9;	// matmul/matmul-hw.mlir:19667:22
  wire [31:0]     b_i_k_7_i_j_9;	// matmul/matmul-hw.mlir:19670:22
  wire [31:0]     c_prev_i_k_7_i_j_9;	// matmul/matmul-hw.mlir:19673:27
  wire            tk_i_k_7_i_j_9;	// matmul/matmul-hw.mlir:19676:23
  wire [31:0]     c_i_k_7_i_j_9;	// matmul/matmul-hw.mlir:19680:22
  reg  [3:0]      i_k_next_3590;	// matmul/matmul-hw.mlir:19685:22
  wire [31:0]     a_i_k_8_i_j_9;	// matmul/matmul-hw.mlir:19697:22
  wire [31:0]     b_i_k_8_i_j_9;	// matmul/matmul-hw.mlir:19700:22
  wire [31:0]     c_prev_i_k_8_i_j_9;	// matmul/matmul-hw.mlir:19703:27
  wire            tk_i_k_8_i_j_9;	// matmul/matmul-hw.mlir:19706:23
  wire [31:0]     c_i_k_8_i_j_9;	// matmul/matmul-hw.mlir:19710:22
  reg  [3:0]      i_k_next_3593;	// matmul/matmul-hw.mlir:19715:22
  wire [31:0]     a_i_k_9_i_j_9;	// matmul/matmul-hw.mlir:19727:22
  wire [31:0]     b_i_k_9_i_j_9;	// matmul/matmul-hw.mlir:19730:22
  wire [31:0]     c_prev_i_k_9_i_j_9;	// matmul/matmul-hw.mlir:19733:27
  wire            tk_i_k_9_i_j_9;	// matmul/matmul-hw.mlir:19736:23
  wire [31:0]     c_i_k_9_i_j_9;	// matmul/matmul-hw.mlir:19740:22
  reg  [3:0]      i_k_next_3596;	// matmul/matmul-hw.mlir:19745:22
  wire [31:0]     a_i_k_10_i_j_9;	// matmul/matmul-hw.mlir:19757:23
  wire [31:0]     b_i_k_10_i_j_9;	// matmul/matmul-hw.mlir:19760:23
  wire [31:0]     c_prev_i_k_10_i_j_9;	// matmul/matmul-hw.mlir:19763:28
  wire            tk_i_k_10_i_j_9;	// matmul/matmul-hw.mlir:19766:24
  wire [31:0]     c_i_k_10_i_j_9;	// matmul/matmul-hw.mlir:19770:23
  reg  [3:0]      i_k_next_3599;	// matmul/matmul-hw.mlir:19775:22
  wire [31:0]     a_i_k_11_i_j_9;	// matmul/matmul-hw.mlir:19787:23
  wire [31:0]     b_i_k_11_i_j_9;	// matmul/matmul-hw.mlir:19790:23
  wire [31:0]     c_prev_i_k_11_i_j_9;	// matmul/matmul-hw.mlir:19793:28
  wire            tk_i_k_11_i_j_9;	// matmul/matmul-hw.mlir:19796:24
  wire [31:0]     c_i_k_11_i_j_9;	// matmul/matmul-hw.mlir:19800:23
  reg  [3:0]      i_k_next_3602;	// matmul/matmul-hw.mlir:19805:22
  wire [31:0]     a_i_k_12_i_j_9;	// matmul/matmul-hw.mlir:19817:23
  wire [31:0]     b_i_k_12_i_j_9;	// matmul/matmul-hw.mlir:19820:23
  wire [31:0]     c_prev_i_k_12_i_j_9;	// matmul/matmul-hw.mlir:19823:28
  wire            tk_i_k_12_i_j_9;	// matmul/matmul-hw.mlir:19826:24
  wire [31:0]     c_i_k_12_i_j_9;	// matmul/matmul-hw.mlir:19830:23
  reg  [3:0]      i_k_next_3605;	// matmul/matmul-hw.mlir:19835:22
  wire [31:0]     a_i_k_13_i_j_9;	// matmul/matmul-hw.mlir:19847:23
  wire [31:0]     b_i_k_13_i_j_9;	// matmul/matmul-hw.mlir:19850:23
  wire [31:0]     c_prev_i_k_13_i_j_9;	// matmul/matmul-hw.mlir:19853:28
  wire            tk_i_k_13_i_j_9;	// matmul/matmul-hw.mlir:19856:24
  wire [31:0]     c_i_k_13_i_j_9;	// matmul/matmul-hw.mlir:19860:23
  reg  [3:0]      i_k_next_3608;	// matmul/matmul-hw.mlir:19865:22
  wire [31:0]     a_i_k_14_i_j_9;	// matmul/matmul-hw.mlir:19877:23
  wire [31:0]     b_i_k_14_i_j_9;	// matmul/matmul-hw.mlir:19880:23
  wire [31:0]     c_prev_i_k_14_i_j_9;	// matmul/matmul-hw.mlir:19883:28
  wire            tk_i_k_14_i_j_9;	// matmul/matmul-hw.mlir:19886:24
  wire [31:0]     c_i_k_14_i_j_9;	// matmul/matmul-hw.mlir:19890:23
  reg  [3:0]      i_k_next_3611;	// matmul/matmul-hw.mlir:19895:22
  wire [31:0]     a_i_k_15_i_j_9;	// matmul/matmul-hw.mlir:19907:23
  wire [31:0]     b_i_k_15_i_j_9;	// matmul/matmul-hw.mlir:19910:23
  wire [31:0]     c_prev_i_k_15_i_j_9;	// matmul/matmul-hw.mlir:19913:28
  wire            tk_i_k_15_i_j_9;	// matmul/matmul-hw.mlir:19916:24
  wire [31:0]     c_i_k_15_i_j_9;	// matmul/matmul-hw.mlir:19920:23
  reg  [3:0]      i_k_next_3614;	// matmul/matmul-hw.mlir:19925:22
  reg  [3:0][3:0] i_delayed_3616;	// matmul/matmul-hw.mlir:19934:23
  reg  [3:0]      i_j_next_3620;	// matmul/matmul-hw.mlir:19953:22
  wire [31:0]     a_i_k_0_i_j_10;	// matmul/matmul-hw.mlir:20052:23
  wire [31:0]     b_i_k_0_i_j_10;	// matmul/matmul-hw.mlir:20055:23
  wire [31:0]     c_prev_i_k_0_i_j_10;	// matmul/matmul-hw.mlir:20058:28
  wire            tk_i_k_0_i_j_10;	// matmul/matmul-hw.mlir:20061:24
  wire [31:0]     c_i_k_0_i_j_10;	// matmul/matmul-hw.mlir:20065:23
  reg  [3:0]      i_k_next_3640;	// matmul/matmul-hw.mlir:20070:22
  wire [31:0]     a_i_k_1_i_j_10;	// matmul/matmul-hw.mlir:20082:23
  wire [31:0]     b_i_k_1_i_j_10;	// matmul/matmul-hw.mlir:20085:23
  wire [31:0]     c_prev_i_k_1_i_j_10;	// matmul/matmul-hw.mlir:20088:28
  wire            tk_i_k_1_i_j_10;	// matmul/matmul-hw.mlir:20091:24
  wire [31:0]     c_i_k_1_i_j_10;	// matmul/matmul-hw.mlir:20095:23
  reg  [3:0]      i_k_next_3643;	// matmul/matmul-hw.mlir:20100:22
  wire [31:0]     a_i_k_2_i_j_10;	// matmul/matmul-hw.mlir:20112:23
  wire [31:0]     b_i_k_2_i_j_10;	// matmul/matmul-hw.mlir:20115:23
  wire [31:0]     c_prev_i_k_2_i_j_10;	// matmul/matmul-hw.mlir:20118:28
  wire            tk_i_k_2_i_j_10;	// matmul/matmul-hw.mlir:20121:24
  wire [31:0]     c_i_k_2_i_j_10;	// matmul/matmul-hw.mlir:20125:23
  reg  [3:0]      i_k_next_3646;	// matmul/matmul-hw.mlir:20130:22
  wire [31:0]     a_i_k_3_i_j_10;	// matmul/matmul-hw.mlir:20142:23
  wire [31:0]     b_i_k_3_i_j_10;	// matmul/matmul-hw.mlir:20145:23
  wire [31:0]     c_prev_i_k_3_i_j_10;	// matmul/matmul-hw.mlir:20148:28
  wire            tk_i_k_3_i_j_10;	// matmul/matmul-hw.mlir:20151:24
  wire [31:0]     c_i_k_3_i_j_10;	// matmul/matmul-hw.mlir:20155:23
  reg  [3:0]      i_k_next_3649;	// matmul/matmul-hw.mlir:20160:22
  wire [31:0]     a_i_k_4_i_j_10;	// matmul/matmul-hw.mlir:20172:23
  wire [31:0]     b_i_k_4_i_j_10;	// matmul/matmul-hw.mlir:20175:23
  wire [31:0]     c_prev_i_k_4_i_j_10;	// matmul/matmul-hw.mlir:20178:28
  wire            tk_i_k_4_i_j_10;	// matmul/matmul-hw.mlir:20181:24
  wire [31:0]     c_i_k_4_i_j_10;	// matmul/matmul-hw.mlir:20185:23
  reg  [3:0]      i_k_next_3652;	// matmul/matmul-hw.mlir:20190:22
  wire [31:0]     a_i_k_5_i_j_10;	// matmul/matmul-hw.mlir:20202:23
  wire [31:0]     b_i_k_5_i_j_10;	// matmul/matmul-hw.mlir:20205:23
  wire [31:0]     c_prev_i_k_5_i_j_10;	// matmul/matmul-hw.mlir:20208:28
  wire            tk_i_k_5_i_j_10;	// matmul/matmul-hw.mlir:20211:24
  wire [31:0]     c_i_k_5_i_j_10;	// matmul/matmul-hw.mlir:20215:23
  reg  [3:0]      i_k_next_3655;	// matmul/matmul-hw.mlir:20220:22
  wire [31:0]     a_i_k_6_i_j_10;	// matmul/matmul-hw.mlir:20232:23
  wire [31:0]     b_i_k_6_i_j_10;	// matmul/matmul-hw.mlir:20235:23
  wire [31:0]     c_prev_i_k_6_i_j_10;	// matmul/matmul-hw.mlir:20238:28
  wire            tk_i_k_6_i_j_10;	// matmul/matmul-hw.mlir:20241:24
  wire [31:0]     c_i_k_6_i_j_10;	// matmul/matmul-hw.mlir:20245:23
  reg  [3:0]      i_k_next_3658;	// matmul/matmul-hw.mlir:20250:22
  wire [31:0]     a_i_k_7_i_j_10;	// matmul/matmul-hw.mlir:20262:23
  wire [31:0]     b_i_k_7_i_j_10;	// matmul/matmul-hw.mlir:20265:23
  wire [31:0]     c_prev_i_k_7_i_j_10;	// matmul/matmul-hw.mlir:20268:28
  wire            tk_i_k_7_i_j_10;	// matmul/matmul-hw.mlir:20271:24
  wire [31:0]     c_i_k_7_i_j_10;	// matmul/matmul-hw.mlir:20275:23
  reg  [3:0]      i_k_next_3661;	// matmul/matmul-hw.mlir:20280:22
  wire [31:0]     a_i_k_8_i_j_10;	// matmul/matmul-hw.mlir:20292:23
  wire [31:0]     b_i_k_8_i_j_10;	// matmul/matmul-hw.mlir:20295:23
  wire [31:0]     c_prev_i_k_8_i_j_10;	// matmul/matmul-hw.mlir:20298:28
  wire            tk_i_k_8_i_j_10;	// matmul/matmul-hw.mlir:20301:24
  wire [31:0]     c_i_k_8_i_j_10;	// matmul/matmul-hw.mlir:20305:23
  reg  [3:0]      i_k_next_3664;	// matmul/matmul-hw.mlir:20310:22
  wire [31:0]     a_i_k_9_i_j_10;	// matmul/matmul-hw.mlir:20322:23
  wire [31:0]     b_i_k_9_i_j_10;	// matmul/matmul-hw.mlir:20325:23
  wire [31:0]     c_prev_i_k_9_i_j_10;	// matmul/matmul-hw.mlir:20328:28
  wire            tk_i_k_9_i_j_10;	// matmul/matmul-hw.mlir:20331:24
  wire [31:0]     c_i_k_9_i_j_10;	// matmul/matmul-hw.mlir:20335:23
  reg  [3:0]      i_k_next_3667;	// matmul/matmul-hw.mlir:20340:22
  wire [31:0]     a_i_k_10_i_j_10;	// matmul/matmul-hw.mlir:20352:24
  wire [31:0]     b_i_k_10_i_j_10;	// matmul/matmul-hw.mlir:20355:24
  wire [31:0]     c_prev_i_k_10_i_j_10;	// matmul/matmul-hw.mlir:20358:29
  wire            tk_i_k_10_i_j_10;	// matmul/matmul-hw.mlir:20361:25
  wire [31:0]     c_i_k_10_i_j_10;	// matmul/matmul-hw.mlir:20365:24
  reg  [3:0]      i_k_next_3670;	// matmul/matmul-hw.mlir:20370:22
  wire [31:0]     a_i_k_11_i_j_10;	// matmul/matmul-hw.mlir:20382:24
  wire [31:0]     b_i_k_11_i_j_10;	// matmul/matmul-hw.mlir:20385:24
  wire [31:0]     c_prev_i_k_11_i_j_10;	// matmul/matmul-hw.mlir:20388:29
  wire            tk_i_k_11_i_j_10;	// matmul/matmul-hw.mlir:20391:25
  wire [31:0]     c_i_k_11_i_j_10;	// matmul/matmul-hw.mlir:20395:24
  reg  [3:0]      i_k_next_3673;	// matmul/matmul-hw.mlir:20400:22
  wire [31:0]     a_i_k_12_i_j_10;	// matmul/matmul-hw.mlir:20412:24
  wire [31:0]     b_i_k_12_i_j_10;	// matmul/matmul-hw.mlir:20415:24
  wire [31:0]     c_prev_i_k_12_i_j_10;	// matmul/matmul-hw.mlir:20418:29
  wire            tk_i_k_12_i_j_10;	// matmul/matmul-hw.mlir:20421:25
  wire [31:0]     c_i_k_12_i_j_10;	// matmul/matmul-hw.mlir:20425:24
  reg  [3:0]      i_k_next_3676;	// matmul/matmul-hw.mlir:20430:22
  wire [31:0]     a_i_k_13_i_j_10;	// matmul/matmul-hw.mlir:20442:24
  wire [31:0]     b_i_k_13_i_j_10;	// matmul/matmul-hw.mlir:20445:24
  wire [31:0]     c_prev_i_k_13_i_j_10;	// matmul/matmul-hw.mlir:20448:29
  wire            tk_i_k_13_i_j_10;	// matmul/matmul-hw.mlir:20451:25
  wire [31:0]     c_i_k_13_i_j_10;	// matmul/matmul-hw.mlir:20455:24
  reg  [3:0]      i_k_next_3679;	// matmul/matmul-hw.mlir:20460:22
  wire [31:0]     a_i_k_14_i_j_10;	// matmul/matmul-hw.mlir:20472:24
  wire [31:0]     b_i_k_14_i_j_10;	// matmul/matmul-hw.mlir:20475:24
  wire [31:0]     c_prev_i_k_14_i_j_10;	// matmul/matmul-hw.mlir:20478:29
  wire            tk_i_k_14_i_j_10;	// matmul/matmul-hw.mlir:20481:25
  wire [31:0]     c_i_k_14_i_j_10;	// matmul/matmul-hw.mlir:20485:24
  reg  [3:0]      i_k_next_3682;	// matmul/matmul-hw.mlir:20490:22
  wire [31:0]     a_i_k_15_i_j_10;	// matmul/matmul-hw.mlir:20502:24
  wire [31:0]     b_i_k_15_i_j_10;	// matmul/matmul-hw.mlir:20505:24
  wire [31:0]     c_prev_i_k_15_i_j_10;	// matmul/matmul-hw.mlir:20508:29
  wire            tk_i_k_15_i_j_10;	// matmul/matmul-hw.mlir:20511:25
  wire [31:0]     c_i_k_15_i_j_10;	// matmul/matmul-hw.mlir:20515:24
  reg  [3:0]      i_k_next_3685;	// matmul/matmul-hw.mlir:20520:22
  reg  [3:0][3:0] i_delayed_3687;	// matmul/matmul-hw.mlir:20529:23
  reg  [3:0]      i_j_next_3691;	// matmul/matmul-hw.mlir:20548:22
  wire [31:0]     a_i_k_0_i_j_11;	// matmul/matmul-hw.mlir:20647:23
  wire [31:0]     b_i_k_0_i_j_11;	// matmul/matmul-hw.mlir:20650:23
  wire [31:0]     c_prev_i_k_0_i_j_11;	// matmul/matmul-hw.mlir:20653:28
  wire            tk_i_k_0_i_j_11;	// matmul/matmul-hw.mlir:20656:24
  wire [31:0]     c_i_k_0_i_j_11;	// matmul/matmul-hw.mlir:20660:23
  reg  [3:0]      i_k_next_3711;	// matmul/matmul-hw.mlir:20665:22
  wire [31:0]     a_i_k_1_i_j_11;	// matmul/matmul-hw.mlir:20677:23
  wire [31:0]     b_i_k_1_i_j_11;	// matmul/matmul-hw.mlir:20680:23
  wire [31:0]     c_prev_i_k_1_i_j_11;	// matmul/matmul-hw.mlir:20683:28
  wire            tk_i_k_1_i_j_11;	// matmul/matmul-hw.mlir:20686:24
  wire [31:0]     c_i_k_1_i_j_11;	// matmul/matmul-hw.mlir:20690:23
  reg  [3:0]      i_k_next_3714;	// matmul/matmul-hw.mlir:20695:22
  wire [31:0]     a_i_k_2_i_j_11;	// matmul/matmul-hw.mlir:20707:23
  wire [31:0]     b_i_k_2_i_j_11;	// matmul/matmul-hw.mlir:20710:23
  wire [31:0]     c_prev_i_k_2_i_j_11;	// matmul/matmul-hw.mlir:20713:28
  wire            tk_i_k_2_i_j_11;	// matmul/matmul-hw.mlir:20716:24
  wire [31:0]     c_i_k_2_i_j_11;	// matmul/matmul-hw.mlir:20720:23
  reg  [3:0]      i_k_next_3717;	// matmul/matmul-hw.mlir:20725:22
  wire [31:0]     a_i_k_3_i_j_11;	// matmul/matmul-hw.mlir:20737:23
  wire [31:0]     b_i_k_3_i_j_11;	// matmul/matmul-hw.mlir:20740:23
  wire [31:0]     c_prev_i_k_3_i_j_11;	// matmul/matmul-hw.mlir:20743:28
  wire            tk_i_k_3_i_j_11;	// matmul/matmul-hw.mlir:20746:24
  wire [31:0]     c_i_k_3_i_j_11;	// matmul/matmul-hw.mlir:20750:23
  reg  [3:0]      i_k_next_3720;	// matmul/matmul-hw.mlir:20755:22
  wire [31:0]     a_i_k_4_i_j_11;	// matmul/matmul-hw.mlir:20767:23
  wire [31:0]     b_i_k_4_i_j_11;	// matmul/matmul-hw.mlir:20770:23
  wire [31:0]     c_prev_i_k_4_i_j_11;	// matmul/matmul-hw.mlir:20773:28
  wire            tk_i_k_4_i_j_11;	// matmul/matmul-hw.mlir:20776:24
  wire [31:0]     c_i_k_4_i_j_11;	// matmul/matmul-hw.mlir:20780:23
  reg  [3:0]      i_k_next_3723;	// matmul/matmul-hw.mlir:20785:22
  wire [31:0]     a_i_k_5_i_j_11;	// matmul/matmul-hw.mlir:20797:23
  wire [31:0]     b_i_k_5_i_j_11;	// matmul/matmul-hw.mlir:20800:23
  wire [31:0]     c_prev_i_k_5_i_j_11;	// matmul/matmul-hw.mlir:20803:28
  wire            tk_i_k_5_i_j_11;	// matmul/matmul-hw.mlir:20806:24
  wire [31:0]     c_i_k_5_i_j_11;	// matmul/matmul-hw.mlir:20810:23
  reg  [3:0]      i_k_next_3726;	// matmul/matmul-hw.mlir:20815:22
  wire [31:0]     a_i_k_6_i_j_11;	// matmul/matmul-hw.mlir:20827:23
  wire [31:0]     b_i_k_6_i_j_11;	// matmul/matmul-hw.mlir:20830:23
  wire [31:0]     c_prev_i_k_6_i_j_11;	// matmul/matmul-hw.mlir:20833:28
  wire            tk_i_k_6_i_j_11;	// matmul/matmul-hw.mlir:20836:24
  wire [31:0]     c_i_k_6_i_j_11;	// matmul/matmul-hw.mlir:20840:23
  reg  [3:0]      i_k_next_3729;	// matmul/matmul-hw.mlir:20845:22
  wire [31:0]     a_i_k_7_i_j_11;	// matmul/matmul-hw.mlir:20857:23
  wire [31:0]     b_i_k_7_i_j_11;	// matmul/matmul-hw.mlir:20860:23
  wire [31:0]     c_prev_i_k_7_i_j_11;	// matmul/matmul-hw.mlir:20863:28
  wire            tk_i_k_7_i_j_11;	// matmul/matmul-hw.mlir:20866:24
  wire [31:0]     c_i_k_7_i_j_11;	// matmul/matmul-hw.mlir:20870:23
  reg  [3:0]      i_k_next_3732;	// matmul/matmul-hw.mlir:20875:22
  wire [31:0]     a_i_k_8_i_j_11;	// matmul/matmul-hw.mlir:20887:23
  wire [31:0]     b_i_k_8_i_j_11;	// matmul/matmul-hw.mlir:20890:23
  wire [31:0]     c_prev_i_k_8_i_j_11;	// matmul/matmul-hw.mlir:20893:28
  wire            tk_i_k_8_i_j_11;	// matmul/matmul-hw.mlir:20896:24
  wire [31:0]     c_i_k_8_i_j_11;	// matmul/matmul-hw.mlir:20900:23
  reg  [3:0]      i_k_next_3735;	// matmul/matmul-hw.mlir:20905:22
  wire [31:0]     a_i_k_9_i_j_11;	// matmul/matmul-hw.mlir:20917:23
  wire [31:0]     b_i_k_9_i_j_11;	// matmul/matmul-hw.mlir:20920:23
  wire [31:0]     c_prev_i_k_9_i_j_11;	// matmul/matmul-hw.mlir:20923:28
  wire            tk_i_k_9_i_j_11;	// matmul/matmul-hw.mlir:20926:24
  wire [31:0]     c_i_k_9_i_j_11;	// matmul/matmul-hw.mlir:20930:23
  reg  [3:0]      i_k_next_3738;	// matmul/matmul-hw.mlir:20935:22
  wire [31:0]     a_i_k_10_i_j_11;	// matmul/matmul-hw.mlir:20947:24
  wire [31:0]     b_i_k_10_i_j_11;	// matmul/matmul-hw.mlir:20950:24
  wire [31:0]     c_prev_i_k_10_i_j_11;	// matmul/matmul-hw.mlir:20953:29
  wire            tk_i_k_10_i_j_11;	// matmul/matmul-hw.mlir:20956:25
  wire [31:0]     c_i_k_10_i_j_11;	// matmul/matmul-hw.mlir:20960:24
  reg  [3:0]      i_k_next_3741;	// matmul/matmul-hw.mlir:20965:22
  wire [31:0]     a_i_k_11_i_j_11;	// matmul/matmul-hw.mlir:20977:24
  wire [31:0]     b_i_k_11_i_j_11;	// matmul/matmul-hw.mlir:20980:24
  wire [31:0]     c_prev_i_k_11_i_j_11;	// matmul/matmul-hw.mlir:20983:29
  wire            tk_i_k_11_i_j_11;	// matmul/matmul-hw.mlir:20986:25
  wire [31:0]     c_i_k_11_i_j_11;	// matmul/matmul-hw.mlir:20990:24
  reg  [3:0]      i_k_next_3744;	// matmul/matmul-hw.mlir:20995:22
  wire [31:0]     a_i_k_12_i_j_11;	// matmul/matmul-hw.mlir:21007:24
  wire [31:0]     b_i_k_12_i_j_11;	// matmul/matmul-hw.mlir:21010:24
  wire [31:0]     c_prev_i_k_12_i_j_11;	// matmul/matmul-hw.mlir:21013:29
  wire            tk_i_k_12_i_j_11;	// matmul/matmul-hw.mlir:21016:25
  wire [31:0]     c_i_k_12_i_j_11;	// matmul/matmul-hw.mlir:21020:24
  reg  [3:0]      i_k_next_3747;	// matmul/matmul-hw.mlir:21025:22
  wire [31:0]     a_i_k_13_i_j_11;	// matmul/matmul-hw.mlir:21037:24
  wire [31:0]     b_i_k_13_i_j_11;	// matmul/matmul-hw.mlir:21040:24
  wire [31:0]     c_prev_i_k_13_i_j_11;	// matmul/matmul-hw.mlir:21043:29
  wire            tk_i_k_13_i_j_11;	// matmul/matmul-hw.mlir:21046:25
  wire [31:0]     c_i_k_13_i_j_11;	// matmul/matmul-hw.mlir:21050:24
  reg  [3:0]      i_k_next_3750;	// matmul/matmul-hw.mlir:21055:22
  wire [31:0]     a_i_k_14_i_j_11;	// matmul/matmul-hw.mlir:21067:24
  wire [31:0]     b_i_k_14_i_j_11;	// matmul/matmul-hw.mlir:21070:24
  wire [31:0]     c_prev_i_k_14_i_j_11;	// matmul/matmul-hw.mlir:21073:29
  wire            tk_i_k_14_i_j_11;	// matmul/matmul-hw.mlir:21076:25
  wire [31:0]     c_i_k_14_i_j_11;	// matmul/matmul-hw.mlir:21080:24
  reg  [3:0]      i_k_next_3753;	// matmul/matmul-hw.mlir:21085:22
  wire [31:0]     a_i_k_15_i_j_11;	// matmul/matmul-hw.mlir:21097:24
  wire [31:0]     b_i_k_15_i_j_11;	// matmul/matmul-hw.mlir:21100:24
  wire [31:0]     c_prev_i_k_15_i_j_11;	// matmul/matmul-hw.mlir:21103:29
  wire            tk_i_k_15_i_j_11;	// matmul/matmul-hw.mlir:21106:25
  wire [31:0]     c_i_k_15_i_j_11;	// matmul/matmul-hw.mlir:21110:24
  reg  [3:0]      i_k_next_3756;	// matmul/matmul-hw.mlir:21115:22
  reg  [3:0][3:0] i_delayed_3758;	// matmul/matmul-hw.mlir:21124:23
  reg  [3:0]      i_j_next_3762;	// matmul/matmul-hw.mlir:21143:22
  wire [31:0]     a_i_k_0_i_j_12;	// matmul/matmul-hw.mlir:21242:23
  wire [31:0]     b_i_k_0_i_j_12;	// matmul/matmul-hw.mlir:21245:23
  wire [31:0]     c_prev_i_k_0_i_j_12;	// matmul/matmul-hw.mlir:21248:28
  wire            tk_i_k_0_i_j_12;	// matmul/matmul-hw.mlir:21251:24
  wire [31:0]     c_i_k_0_i_j_12;	// matmul/matmul-hw.mlir:21255:23
  reg  [3:0]      i_k_next_3782;	// matmul/matmul-hw.mlir:21260:22
  wire [31:0]     a_i_k_1_i_j_12;	// matmul/matmul-hw.mlir:21272:23
  wire [31:0]     b_i_k_1_i_j_12;	// matmul/matmul-hw.mlir:21275:23
  wire [31:0]     c_prev_i_k_1_i_j_12;	// matmul/matmul-hw.mlir:21278:28
  wire            tk_i_k_1_i_j_12;	// matmul/matmul-hw.mlir:21281:24
  wire [31:0]     c_i_k_1_i_j_12;	// matmul/matmul-hw.mlir:21285:23
  reg  [3:0]      i_k_next_3785;	// matmul/matmul-hw.mlir:21290:22
  wire [31:0]     a_i_k_2_i_j_12;	// matmul/matmul-hw.mlir:21302:23
  wire [31:0]     b_i_k_2_i_j_12;	// matmul/matmul-hw.mlir:21305:23
  wire [31:0]     c_prev_i_k_2_i_j_12;	// matmul/matmul-hw.mlir:21308:28
  wire            tk_i_k_2_i_j_12;	// matmul/matmul-hw.mlir:21311:24
  wire [31:0]     c_i_k_2_i_j_12;	// matmul/matmul-hw.mlir:21315:23
  reg  [3:0]      i_k_next_3788;	// matmul/matmul-hw.mlir:21320:22
  wire [31:0]     a_i_k_3_i_j_12;	// matmul/matmul-hw.mlir:21332:23
  wire [31:0]     b_i_k_3_i_j_12;	// matmul/matmul-hw.mlir:21335:23
  wire [31:0]     c_prev_i_k_3_i_j_12;	// matmul/matmul-hw.mlir:21338:28
  wire            tk_i_k_3_i_j_12;	// matmul/matmul-hw.mlir:21341:24
  wire [31:0]     c_i_k_3_i_j_12;	// matmul/matmul-hw.mlir:21345:23
  reg  [3:0]      i_k_next_3791;	// matmul/matmul-hw.mlir:21350:22
  wire [31:0]     a_i_k_4_i_j_12;	// matmul/matmul-hw.mlir:21362:23
  wire [31:0]     b_i_k_4_i_j_12;	// matmul/matmul-hw.mlir:21365:23
  wire [31:0]     c_prev_i_k_4_i_j_12;	// matmul/matmul-hw.mlir:21368:28
  wire            tk_i_k_4_i_j_12;	// matmul/matmul-hw.mlir:21371:24
  wire [31:0]     c_i_k_4_i_j_12;	// matmul/matmul-hw.mlir:21375:23
  reg  [3:0]      i_k_next_3794;	// matmul/matmul-hw.mlir:21380:22
  wire [31:0]     a_i_k_5_i_j_12;	// matmul/matmul-hw.mlir:21392:23
  wire [31:0]     b_i_k_5_i_j_12;	// matmul/matmul-hw.mlir:21395:23
  wire [31:0]     c_prev_i_k_5_i_j_12;	// matmul/matmul-hw.mlir:21398:28
  wire            tk_i_k_5_i_j_12;	// matmul/matmul-hw.mlir:21401:24
  wire [31:0]     c_i_k_5_i_j_12;	// matmul/matmul-hw.mlir:21405:23
  reg  [3:0]      i_k_next_3797;	// matmul/matmul-hw.mlir:21410:22
  wire [31:0]     a_i_k_6_i_j_12;	// matmul/matmul-hw.mlir:21422:23
  wire [31:0]     b_i_k_6_i_j_12;	// matmul/matmul-hw.mlir:21425:23
  wire [31:0]     c_prev_i_k_6_i_j_12;	// matmul/matmul-hw.mlir:21428:28
  wire            tk_i_k_6_i_j_12;	// matmul/matmul-hw.mlir:21431:24
  wire [31:0]     c_i_k_6_i_j_12;	// matmul/matmul-hw.mlir:21435:23
  reg  [3:0]      i_k_next_3800;	// matmul/matmul-hw.mlir:21440:22
  wire [31:0]     a_i_k_7_i_j_12;	// matmul/matmul-hw.mlir:21452:23
  wire [31:0]     b_i_k_7_i_j_12;	// matmul/matmul-hw.mlir:21455:23
  wire [31:0]     c_prev_i_k_7_i_j_12;	// matmul/matmul-hw.mlir:21458:28
  wire            tk_i_k_7_i_j_12;	// matmul/matmul-hw.mlir:21461:24
  wire [31:0]     c_i_k_7_i_j_12;	// matmul/matmul-hw.mlir:21465:23
  reg  [3:0]      i_k_next_3803;	// matmul/matmul-hw.mlir:21470:22
  wire [31:0]     a_i_k_8_i_j_12;	// matmul/matmul-hw.mlir:21482:23
  wire [31:0]     b_i_k_8_i_j_12;	// matmul/matmul-hw.mlir:21485:23
  wire [31:0]     c_prev_i_k_8_i_j_12;	// matmul/matmul-hw.mlir:21488:28
  wire            tk_i_k_8_i_j_12;	// matmul/matmul-hw.mlir:21491:24
  wire [31:0]     c_i_k_8_i_j_12;	// matmul/matmul-hw.mlir:21495:23
  reg  [3:0]      i_k_next_3806;	// matmul/matmul-hw.mlir:21500:22
  wire [31:0]     a_i_k_9_i_j_12;	// matmul/matmul-hw.mlir:21512:23
  wire [31:0]     b_i_k_9_i_j_12;	// matmul/matmul-hw.mlir:21515:23
  wire [31:0]     c_prev_i_k_9_i_j_12;	// matmul/matmul-hw.mlir:21518:28
  wire            tk_i_k_9_i_j_12;	// matmul/matmul-hw.mlir:21521:24
  wire [31:0]     c_i_k_9_i_j_12;	// matmul/matmul-hw.mlir:21525:23
  reg  [3:0]      i_k_next_3809;	// matmul/matmul-hw.mlir:21530:22
  wire [31:0]     a_i_k_10_i_j_12;	// matmul/matmul-hw.mlir:21542:24
  wire [31:0]     b_i_k_10_i_j_12;	// matmul/matmul-hw.mlir:21545:24
  wire [31:0]     c_prev_i_k_10_i_j_12;	// matmul/matmul-hw.mlir:21548:29
  wire            tk_i_k_10_i_j_12;	// matmul/matmul-hw.mlir:21551:25
  wire [31:0]     c_i_k_10_i_j_12;	// matmul/matmul-hw.mlir:21555:24
  reg  [3:0]      i_k_next_3812;	// matmul/matmul-hw.mlir:21560:22
  wire [31:0]     a_i_k_11_i_j_12;	// matmul/matmul-hw.mlir:21572:24
  wire [31:0]     b_i_k_11_i_j_12;	// matmul/matmul-hw.mlir:21575:24
  wire [31:0]     c_prev_i_k_11_i_j_12;	// matmul/matmul-hw.mlir:21578:29
  wire            tk_i_k_11_i_j_12;	// matmul/matmul-hw.mlir:21581:25
  wire [31:0]     c_i_k_11_i_j_12;	// matmul/matmul-hw.mlir:21585:24
  reg  [3:0]      i_k_next_3815;	// matmul/matmul-hw.mlir:21590:22
  wire [31:0]     a_i_k_12_i_j_12;	// matmul/matmul-hw.mlir:21602:24
  wire [31:0]     b_i_k_12_i_j_12;	// matmul/matmul-hw.mlir:21605:24
  wire [31:0]     c_prev_i_k_12_i_j_12;	// matmul/matmul-hw.mlir:21608:29
  wire            tk_i_k_12_i_j_12;	// matmul/matmul-hw.mlir:21611:25
  wire [31:0]     c_i_k_12_i_j_12;	// matmul/matmul-hw.mlir:21615:24
  reg  [3:0]      i_k_next_3818;	// matmul/matmul-hw.mlir:21620:22
  wire [31:0]     a_i_k_13_i_j_12;	// matmul/matmul-hw.mlir:21632:24
  wire [31:0]     b_i_k_13_i_j_12;	// matmul/matmul-hw.mlir:21635:24
  wire [31:0]     c_prev_i_k_13_i_j_12;	// matmul/matmul-hw.mlir:21638:29
  wire            tk_i_k_13_i_j_12;	// matmul/matmul-hw.mlir:21641:25
  wire [31:0]     c_i_k_13_i_j_12;	// matmul/matmul-hw.mlir:21645:24
  reg  [3:0]      i_k_next_3821;	// matmul/matmul-hw.mlir:21650:22
  wire [31:0]     a_i_k_14_i_j_12;	// matmul/matmul-hw.mlir:21662:24
  wire [31:0]     b_i_k_14_i_j_12;	// matmul/matmul-hw.mlir:21665:24
  wire [31:0]     c_prev_i_k_14_i_j_12;	// matmul/matmul-hw.mlir:21668:29
  wire            tk_i_k_14_i_j_12;	// matmul/matmul-hw.mlir:21671:25
  wire [31:0]     c_i_k_14_i_j_12;	// matmul/matmul-hw.mlir:21675:24
  reg  [3:0]      i_k_next_3824;	// matmul/matmul-hw.mlir:21680:22
  wire [31:0]     a_i_k_15_i_j_12;	// matmul/matmul-hw.mlir:21692:24
  wire [31:0]     b_i_k_15_i_j_12;	// matmul/matmul-hw.mlir:21695:24
  wire [31:0]     c_prev_i_k_15_i_j_12;	// matmul/matmul-hw.mlir:21698:29
  wire            tk_i_k_15_i_j_12;	// matmul/matmul-hw.mlir:21701:25
  wire [31:0]     c_i_k_15_i_j_12;	// matmul/matmul-hw.mlir:21705:24
  reg  [3:0]      i_k_next_3827;	// matmul/matmul-hw.mlir:21710:22
  reg  [31:0]     _T_3829;	// matmul/matmul-hw.mlir:21718:13
  reg  [3:0][3:0] i_delayed_3834;	// matmul/matmul-hw.mlir:21734:23
  reg  [3:0]      i_j_next_3838;	// matmul/matmul-hw.mlir:21753:22
  wire [31:0]     a_i_k_0_i_j_13;	// matmul/matmul-hw.mlir:21852:23
  wire [31:0]     b_i_k_0_i_j_13;	// matmul/matmul-hw.mlir:21855:23
  wire [31:0]     c_prev_i_k_0_i_j_13;	// matmul/matmul-hw.mlir:21858:28
  wire            tk_i_k_0_i_j_13;	// matmul/matmul-hw.mlir:21861:24
  wire [31:0]     c_i_k_0_i_j_13;	// matmul/matmul-hw.mlir:21865:23
  reg  [3:0]      i_k_next_3858;	// matmul/matmul-hw.mlir:21870:22
  wire [31:0]     a_i_k_1_i_j_13;	// matmul/matmul-hw.mlir:21882:23
  wire [31:0]     b_i_k_1_i_j_13;	// matmul/matmul-hw.mlir:21885:23
  wire [31:0]     c_prev_i_k_1_i_j_13;	// matmul/matmul-hw.mlir:21888:28
  wire            tk_i_k_1_i_j_13;	// matmul/matmul-hw.mlir:21891:24
  wire [31:0]     c_i_k_1_i_j_13;	// matmul/matmul-hw.mlir:21895:23
  reg  [3:0]      i_k_next_3861;	// matmul/matmul-hw.mlir:21900:22
  wire [31:0]     a_i_k_2_i_j_13;	// matmul/matmul-hw.mlir:21912:23
  wire [31:0]     b_i_k_2_i_j_13;	// matmul/matmul-hw.mlir:21915:23
  wire [31:0]     c_prev_i_k_2_i_j_13;	// matmul/matmul-hw.mlir:21918:28
  wire            tk_i_k_2_i_j_13;	// matmul/matmul-hw.mlir:21921:24
  wire [31:0]     c_i_k_2_i_j_13;	// matmul/matmul-hw.mlir:21925:23
  reg  [3:0]      i_k_next_3864;	// matmul/matmul-hw.mlir:21930:22
  wire [31:0]     a_i_k_3_i_j_13;	// matmul/matmul-hw.mlir:21942:23
  wire [31:0]     b_i_k_3_i_j_13;	// matmul/matmul-hw.mlir:21945:23
  wire [31:0]     c_prev_i_k_3_i_j_13;	// matmul/matmul-hw.mlir:21948:28
  wire            tk_i_k_3_i_j_13;	// matmul/matmul-hw.mlir:21951:24
  wire [31:0]     c_i_k_3_i_j_13;	// matmul/matmul-hw.mlir:21955:23
  reg  [3:0]      i_k_next_3867;	// matmul/matmul-hw.mlir:21960:22
  wire [31:0]     a_i_k_4_i_j_13;	// matmul/matmul-hw.mlir:21972:23
  wire [31:0]     b_i_k_4_i_j_13;	// matmul/matmul-hw.mlir:21975:23
  wire [31:0]     c_prev_i_k_4_i_j_13;	// matmul/matmul-hw.mlir:21978:28
  wire            tk_i_k_4_i_j_13;	// matmul/matmul-hw.mlir:21981:24
  wire [31:0]     c_i_k_4_i_j_13;	// matmul/matmul-hw.mlir:21985:23
  reg  [3:0]      i_k_next_3870;	// matmul/matmul-hw.mlir:21990:22
  wire [31:0]     a_i_k_5_i_j_13;	// matmul/matmul-hw.mlir:22002:23
  wire [31:0]     b_i_k_5_i_j_13;	// matmul/matmul-hw.mlir:22005:23
  wire [31:0]     c_prev_i_k_5_i_j_13;	// matmul/matmul-hw.mlir:22008:28
  wire            tk_i_k_5_i_j_13;	// matmul/matmul-hw.mlir:22011:24
  wire [31:0]     c_i_k_5_i_j_13;	// matmul/matmul-hw.mlir:22015:23
  reg  [3:0]      i_k_next_3873;	// matmul/matmul-hw.mlir:22020:22
  wire [31:0]     a_i_k_6_i_j_13;	// matmul/matmul-hw.mlir:22032:23
  wire [31:0]     b_i_k_6_i_j_13;	// matmul/matmul-hw.mlir:22035:23
  wire [31:0]     c_prev_i_k_6_i_j_13;	// matmul/matmul-hw.mlir:22038:28
  wire            tk_i_k_6_i_j_13;	// matmul/matmul-hw.mlir:22041:24
  wire [31:0]     c_i_k_6_i_j_13;	// matmul/matmul-hw.mlir:22045:23
  reg  [3:0]      i_k_next_3876;	// matmul/matmul-hw.mlir:22050:22
  wire [31:0]     a_i_k_7_i_j_13;	// matmul/matmul-hw.mlir:22062:23
  wire [31:0]     b_i_k_7_i_j_13;	// matmul/matmul-hw.mlir:22065:23
  wire [31:0]     c_prev_i_k_7_i_j_13;	// matmul/matmul-hw.mlir:22068:28
  wire            tk_i_k_7_i_j_13;	// matmul/matmul-hw.mlir:22071:24
  wire [31:0]     c_i_k_7_i_j_13;	// matmul/matmul-hw.mlir:22075:23
  reg  [3:0]      i_k_next_3879;	// matmul/matmul-hw.mlir:22080:22
  wire [31:0]     a_i_k_8_i_j_13;	// matmul/matmul-hw.mlir:22092:23
  wire [31:0]     b_i_k_8_i_j_13;	// matmul/matmul-hw.mlir:22095:23
  wire [31:0]     c_prev_i_k_8_i_j_13;	// matmul/matmul-hw.mlir:22098:28
  wire            tk_i_k_8_i_j_13;	// matmul/matmul-hw.mlir:22101:24
  wire [31:0]     c_i_k_8_i_j_13;	// matmul/matmul-hw.mlir:22105:23
  reg  [3:0]      i_k_next_3882;	// matmul/matmul-hw.mlir:22110:22
  wire [31:0]     a_i_k_9_i_j_13;	// matmul/matmul-hw.mlir:22122:23
  wire [31:0]     b_i_k_9_i_j_13;	// matmul/matmul-hw.mlir:22125:23
  wire [31:0]     c_prev_i_k_9_i_j_13;	// matmul/matmul-hw.mlir:22128:28
  wire            tk_i_k_9_i_j_13;	// matmul/matmul-hw.mlir:22131:24
  wire [31:0]     c_i_k_9_i_j_13;	// matmul/matmul-hw.mlir:22135:23
  reg  [3:0]      i_k_next_3885;	// matmul/matmul-hw.mlir:22140:22
  wire [31:0]     a_i_k_10_i_j_13;	// matmul/matmul-hw.mlir:22152:24
  wire [31:0]     b_i_k_10_i_j_13;	// matmul/matmul-hw.mlir:22155:24
  wire [31:0]     c_prev_i_k_10_i_j_13;	// matmul/matmul-hw.mlir:22158:29
  wire            tk_i_k_10_i_j_13;	// matmul/matmul-hw.mlir:22161:25
  wire [31:0]     c_i_k_10_i_j_13;	// matmul/matmul-hw.mlir:22165:24
  reg  [3:0]      i_k_next_3888;	// matmul/matmul-hw.mlir:22170:22
  wire [31:0]     a_i_k_11_i_j_13;	// matmul/matmul-hw.mlir:22182:24
  wire [31:0]     b_i_k_11_i_j_13;	// matmul/matmul-hw.mlir:22185:24
  wire [31:0]     c_prev_i_k_11_i_j_13;	// matmul/matmul-hw.mlir:22188:29
  wire            tk_i_k_11_i_j_13;	// matmul/matmul-hw.mlir:22191:25
  wire [31:0]     c_i_k_11_i_j_13;	// matmul/matmul-hw.mlir:22195:24
  reg  [3:0]      i_k_next_3891;	// matmul/matmul-hw.mlir:22200:22
  wire [31:0]     a_i_k_12_i_j_13;	// matmul/matmul-hw.mlir:22212:24
  wire [31:0]     b_i_k_12_i_j_13;	// matmul/matmul-hw.mlir:22215:24
  wire [31:0]     c_prev_i_k_12_i_j_13;	// matmul/matmul-hw.mlir:22218:29
  wire            tk_i_k_12_i_j_13;	// matmul/matmul-hw.mlir:22221:25
  wire [31:0]     c_i_k_12_i_j_13;	// matmul/matmul-hw.mlir:22225:24
  reg  [3:0]      i_k_next_3894;	// matmul/matmul-hw.mlir:22230:22
  wire [31:0]     a_i_k_13_i_j_13;	// matmul/matmul-hw.mlir:22242:24
  wire [31:0]     b_i_k_13_i_j_13;	// matmul/matmul-hw.mlir:22245:24
  wire [31:0]     c_prev_i_k_13_i_j_13;	// matmul/matmul-hw.mlir:22248:29
  wire            tk_i_k_13_i_j_13;	// matmul/matmul-hw.mlir:22251:25
  wire [31:0]     c_i_k_13_i_j_13;	// matmul/matmul-hw.mlir:22255:24
  reg  [3:0]      i_k_next_3897;	// matmul/matmul-hw.mlir:22260:22
  wire [31:0]     a_i_k_14_i_j_13;	// matmul/matmul-hw.mlir:22272:24
  wire [31:0]     b_i_k_14_i_j_13;	// matmul/matmul-hw.mlir:22275:24
  wire [31:0]     c_prev_i_k_14_i_j_13;	// matmul/matmul-hw.mlir:22278:29
  wire            tk_i_k_14_i_j_13;	// matmul/matmul-hw.mlir:22281:25
  wire [31:0]     c_i_k_14_i_j_13;	// matmul/matmul-hw.mlir:22285:24
  reg  [3:0]      i_k_next_3900;	// matmul/matmul-hw.mlir:22290:22
  wire [31:0]     a_i_k_15_i_j_13;	// matmul/matmul-hw.mlir:22302:24
  wire [31:0]     b_i_k_15_i_j_13;	// matmul/matmul-hw.mlir:22305:24
  wire [31:0]     c_prev_i_k_15_i_j_13;	// matmul/matmul-hw.mlir:22308:29
  wire            tk_i_k_15_i_j_13;	// matmul/matmul-hw.mlir:22311:25
  wire [31:0]     c_i_k_15_i_j_13;	// matmul/matmul-hw.mlir:22315:24
  reg  [3:0]      i_k_next_3903;	// matmul/matmul-hw.mlir:22320:22
  reg  [32:0]     _T_3905;	// matmul/matmul-hw.mlir:22328:13
  reg  [3:0][3:0] i_delayed_3910;	// matmul/matmul-hw.mlir:22344:23
  reg  [3:0]      i_j_next_3914;	// matmul/matmul-hw.mlir:22363:22
  wire [31:0]     a_i_k_0_i_j_14;	// matmul/matmul-hw.mlir:22462:23
  wire [31:0]     b_i_k_0_i_j_14;	// matmul/matmul-hw.mlir:22465:23
  wire [31:0]     c_prev_i_k_0_i_j_14;	// matmul/matmul-hw.mlir:22468:28
  wire            tk_i_k_0_i_j_14;	// matmul/matmul-hw.mlir:22471:24
  wire [31:0]     c_i_k_0_i_j_14;	// matmul/matmul-hw.mlir:22475:23
  reg  [3:0]      i_k_next_3934;	// matmul/matmul-hw.mlir:22480:22
  wire [31:0]     a_i_k_1_i_j_14;	// matmul/matmul-hw.mlir:22492:23
  wire [31:0]     b_i_k_1_i_j_14;	// matmul/matmul-hw.mlir:22495:23
  wire [31:0]     c_prev_i_k_1_i_j_14;	// matmul/matmul-hw.mlir:22498:28
  wire            tk_i_k_1_i_j_14;	// matmul/matmul-hw.mlir:22501:24
  wire [31:0]     c_i_k_1_i_j_14;	// matmul/matmul-hw.mlir:22505:23
  reg  [3:0]      i_k_next_3937;	// matmul/matmul-hw.mlir:22510:22
  wire [31:0]     a_i_k_2_i_j_14;	// matmul/matmul-hw.mlir:22522:23
  wire [31:0]     b_i_k_2_i_j_14;	// matmul/matmul-hw.mlir:22525:23
  wire [31:0]     c_prev_i_k_2_i_j_14;	// matmul/matmul-hw.mlir:22528:28
  wire            tk_i_k_2_i_j_14;	// matmul/matmul-hw.mlir:22531:24
  wire [31:0]     c_i_k_2_i_j_14;	// matmul/matmul-hw.mlir:22535:23
  reg  [3:0]      i_k_next_3940;	// matmul/matmul-hw.mlir:22540:22
  wire [31:0]     a_i_k_3_i_j_14;	// matmul/matmul-hw.mlir:22552:23
  wire [31:0]     b_i_k_3_i_j_14;	// matmul/matmul-hw.mlir:22555:23
  wire [31:0]     c_prev_i_k_3_i_j_14;	// matmul/matmul-hw.mlir:22558:28
  wire            tk_i_k_3_i_j_14;	// matmul/matmul-hw.mlir:22561:24
  wire [31:0]     c_i_k_3_i_j_14;	// matmul/matmul-hw.mlir:22565:23
  reg  [3:0]      i_k_next_3943;	// matmul/matmul-hw.mlir:22570:22
  wire [31:0]     a_i_k_4_i_j_14;	// matmul/matmul-hw.mlir:22582:23
  wire [31:0]     b_i_k_4_i_j_14;	// matmul/matmul-hw.mlir:22585:23
  wire [31:0]     c_prev_i_k_4_i_j_14;	// matmul/matmul-hw.mlir:22588:28
  wire            tk_i_k_4_i_j_14;	// matmul/matmul-hw.mlir:22591:24
  wire [31:0]     c_i_k_4_i_j_14;	// matmul/matmul-hw.mlir:22595:23
  reg  [3:0]      i_k_next_3946;	// matmul/matmul-hw.mlir:22600:22
  wire [31:0]     a_i_k_5_i_j_14;	// matmul/matmul-hw.mlir:22612:23
  wire [31:0]     b_i_k_5_i_j_14;	// matmul/matmul-hw.mlir:22615:23
  wire [31:0]     c_prev_i_k_5_i_j_14;	// matmul/matmul-hw.mlir:22618:28
  wire            tk_i_k_5_i_j_14;	// matmul/matmul-hw.mlir:22621:24
  wire [31:0]     c_i_k_5_i_j_14;	// matmul/matmul-hw.mlir:22625:23
  reg  [3:0]      i_k_next_3949;	// matmul/matmul-hw.mlir:22630:22
  wire [31:0]     a_i_k_6_i_j_14;	// matmul/matmul-hw.mlir:22642:23
  wire [31:0]     b_i_k_6_i_j_14;	// matmul/matmul-hw.mlir:22645:23
  wire [31:0]     c_prev_i_k_6_i_j_14;	// matmul/matmul-hw.mlir:22648:28
  wire            tk_i_k_6_i_j_14;	// matmul/matmul-hw.mlir:22651:24
  wire [31:0]     c_i_k_6_i_j_14;	// matmul/matmul-hw.mlir:22655:23
  reg  [3:0]      i_k_next_3952;	// matmul/matmul-hw.mlir:22660:22
  wire [31:0]     a_i_k_7_i_j_14;	// matmul/matmul-hw.mlir:22672:23
  wire [31:0]     b_i_k_7_i_j_14;	// matmul/matmul-hw.mlir:22675:23
  wire [31:0]     c_prev_i_k_7_i_j_14;	// matmul/matmul-hw.mlir:22678:28
  wire            tk_i_k_7_i_j_14;	// matmul/matmul-hw.mlir:22681:24
  wire [31:0]     c_i_k_7_i_j_14;	// matmul/matmul-hw.mlir:22685:23
  reg  [3:0]      i_k_next_3955;	// matmul/matmul-hw.mlir:22690:22
  wire [31:0]     a_i_k_8_i_j_14;	// matmul/matmul-hw.mlir:22702:23
  wire [31:0]     b_i_k_8_i_j_14;	// matmul/matmul-hw.mlir:22705:23
  wire [31:0]     c_prev_i_k_8_i_j_14;	// matmul/matmul-hw.mlir:22708:28
  wire            tk_i_k_8_i_j_14;	// matmul/matmul-hw.mlir:22711:24
  wire [31:0]     c_i_k_8_i_j_14;	// matmul/matmul-hw.mlir:22715:23
  reg  [3:0]      i_k_next_3958;	// matmul/matmul-hw.mlir:22720:22
  wire [31:0]     a_i_k_9_i_j_14;	// matmul/matmul-hw.mlir:22732:23
  wire [31:0]     b_i_k_9_i_j_14;	// matmul/matmul-hw.mlir:22735:23
  wire [31:0]     c_prev_i_k_9_i_j_14;	// matmul/matmul-hw.mlir:22738:28
  wire            tk_i_k_9_i_j_14;	// matmul/matmul-hw.mlir:22741:24
  wire [31:0]     c_i_k_9_i_j_14;	// matmul/matmul-hw.mlir:22745:23
  reg  [3:0]      i_k_next_3961;	// matmul/matmul-hw.mlir:22750:22
  wire [31:0]     a_i_k_10_i_j_14;	// matmul/matmul-hw.mlir:22762:24
  wire [31:0]     b_i_k_10_i_j_14;	// matmul/matmul-hw.mlir:22765:24
  wire [31:0]     c_prev_i_k_10_i_j_14;	// matmul/matmul-hw.mlir:22768:29
  wire            tk_i_k_10_i_j_14;	// matmul/matmul-hw.mlir:22771:25
  wire [31:0]     c_i_k_10_i_j_14;	// matmul/matmul-hw.mlir:22775:24
  reg  [3:0]      i_k_next_3964;	// matmul/matmul-hw.mlir:22780:22
  wire [31:0]     a_i_k_11_i_j_14;	// matmul/matmul-hw.mlir:22792:24
  wire [31:0]     b_i_k_11_i_j_14;	// matmul/matmul-hw.mlir:22795:24
  wire [31:0]     c_prev_i_k_11_i_j_14;	// matmul/matmul-hw.mlir:22798:29
  wire            tk_i_k_11_i_j_14;	// matmul/matmul-hw.mlir:22801:25
  wire [31:0]     c_i_k_11_i_j_14;	// matmul/matmul-hw.mlir:22805:24
  reg  [3:0]      i_k_next_3967;	// matmul/matmul-hw.mlir:22810:22
  wire [31:0]     a_i_k_12_i_j_14;	// matmul/matmul-hw.mlir:22822:24
  wire [31:0]     b_i_k_12_i_j_14;	// matmul/matmul-hw.mlir:22825:24
  wire [31:0]     c_prev_i_k_12_i_j_14;	// matmul/matmul-hw.mlir:22828:29
  wire            tk_i_k_12_i_j_14;	// matmul/matmul-hw.mlir:22831:25
  wire [31:0]     c_i_k_12_i_j_14;	// matmul/matmul-hw.mlir:22835:24
  reg  [3:0]      i_k_next_3970;	// matmul/matmul-hw.mlir:22840:22
  wire [31:0]     a_i_k_13_i_j_14;	// matmul/matmul-hw.mlir:22852:24
  wire [31:0]     b_i_k_13_i_j_14;	// matmul/matmul-hw.mlir:22855:24
  wire [31:0]     c_prev_i_k_13_i_j_14;	// matmul/matmul-hw.mlir:22858:29
  wire            tk_i_k_13_i_j_14;	// matmul/matmul-hw.mlir:22861:25
  wire [31:0]     c_i_k_13_i_j_14;	// matmul/matmul-hw.mlir:22865:24
  reg  [3:0]      i_k_next_3973;	// matmul/matmul-hw.mlir:22870:22
  wire [31:0]     a_i_k_14_i_j_14;	// matmul/matmul-hw.mlir:22882:24
  wire [31:0]     b_i_k_14_i_j_14;	// matmul/matmul-hw.mlir:22885:24
  wire [31:0]     c_prev_i_k_14_i_j_14;	// matmul/matmul-hw.mlir:22888:29
  wire            tk_i_k_14_i_j_14;	// matmul/matmul-hw.mlir:22891:25
  wire [31:0]     c_i_k_14_i_j_14;	// matmul/matmul-hw.mlir:22895:24
  reg  [3:0]      i_k_next_3976;	// matmul/matmul-hw.mlir:22900:22
  wire [31:0]     a_i_k_15_i_j_14;	// matmul/matmul-hw.mlir:22912:24
  wire [31:0]     b_i_k_15_i_j_14;	// matmul/matmul-hw.mlir:22915:24
  wire [31:0]     c_prev_i_k_15_i_j_14;	// matmul/matmul-hw.mlir:22918:29
  wire            tk_i_k_15_i_j_14;	// matmul/matmul-hw.mlir:22921:25
  wire [31:0]     c_i_k_15_i_j_14;	// matmul/matmul-hw.mlir:22925:24
  reg  [3:0]      i_k_next_3979;	// matmul/matmul-hw.mlir:22930:22
  reg  [33:0]     _T_3981;	// matmul/matmul-hw.mlir:22938:13
  reg  [3:0][3:0] i_delayed_3986;	// matmul/matmul-hw.mlir:22954:23
  reg  [3:0]      i_j_next_3990;	// matmul/matmul-hw.mlir:22973:22
  wire [31:0]     a_i_k_0_i_j_15;	// matmul/matmul-hw.mlir:23072:23
  wire [31:0]     b_i_k_0_i_j_15;	// matmul/matmul-hw.mlir:23075:23
  wire [31:0]     c_prev_i_k_0_i_j_15;	// matmul/matmul-hw.mlir:23078:28
  wire            tk_i_k_0_i_j_15;	// matmul/matmul-hw.mlir:23081:24
  wire [31:0]     c_i_k_0_i_j_15;	// matmul/matmul-hw.mlir:23085:23
  reg  [3:0]      i_k_next_4010;	// matmul/matmul-hw.mlir:23090:22
  wire [31:0]     a_i_k_1_i_j_15;	// matmul/matmul-hw.mlir:23102:23
  wire [31:0]     b_i_k_1_i_j_15;	// matmul/matmul-hw.mlir:23105:23
  wire [31:0]     c_prev_i_k_1_i_j_15;	// matmul/matmul-hw.mlir:23108:28
  wire            tk_i_k_1_i_j_15;	// matmul/matmul-hw.mlir:23111:24
  wire [31:0]     c_i_k_1_i_j_15;	// matmul/matmul-hw.mlir:23115:23
  reg  [3:0]      i_k_next_4013;	// matmul/matmul-hw.mlir:23120:22
  wire [31:0]     a_i_k_2_i_j_15;	// matmul/matmul-hw.mlir:23132:23
  wire [31:0]     b_i_k_2_i_j_15;	// matmul/matmul-hw.mlir:23135:23
  wire [31:0]     c_prev_i_k_2_i_j_15;	// matmul/matmul-hw.mlir:23138:28
  wire            tk_i_k_2_i_j_15;	// matmul/matmul-hw.mlir:23141:24
  wire [31:0]     c_i_k_2_i_j_15;	// matmul/matmul-hw.mlir:23145:23
  reg  [3:0]      i_k_next_4016;	// matmul/matmul-hw.mlir:23150:22
  wire [31:0]     a_i_k_3_i_j_15;	// matmul/matmul-hw.mlir:23162:23
  wire [31:0]     b_i_k_3_i_j_15;	// matmul/matmul-hw.mlir:23165:23
  wire [31:0]     c_prev_i_k_3_i_j_15;	// matmul/matmul-hw.mlir:23168:28
  wire            tk_i_k_3_i_j_15;	// matmul/matmul-hw.mlir:23171:24
  wire [31:0]     c_i_k_3_i_j_15;	// matmul/matmul-hw.mlir:23175:23
  reg  [3:0]      i_k_next_4019;	// matmul/matmul-hw.mlir:23180:22
  wire [31:0]     a_i_k_4_i_j_15;	// matmul/matmul-hw.mlir:23192:23
  wire [31:0]     b_i_k_4_i_j_15;	// matmul/matmul-hw.mlir:23195:23
  wire [31:0]     c_prev_i_k_4_i_j_15;	// matmul/matmul-hw.mlir:23198:28
  wire            tk_i_k_4_i_j_15;	// matmul/matmul-hw.mlir:23201:24
  wire [31:0]     c_i_k_4_i_j_15;	// matmul/matmul-hw.mlir:23205:23
  reg  [3:0]      i_k_next_4022;	// matmul/matmul-hw.mlir:23210:22
  wire [31:0]     a_i_k_5_i_j_15;	// matmul/matmul-hw.mlir:23222:23
  wire [31:0]     b_i_k_5_i_j_15;	// matmul/matmul-hw.mlir:23225:23
  wire [31:0]     c_prev_i_k_5_i_j_15;	// matmul/matmul-hw.mlir:23228:28
  wire            tk_i_k_5_i_j_15;	// matmul/matmul-hw.mlir:23231:24
  wire [31:0]     c_i_k_5_i_j_15;	// matmul/matmul-hw.mlir:23235:23
  reg  [3:0]      i_k_next_4025;	// matmul/matmul-hw.mlir:23240:22
  wire [31:0]     a_i_k_6_i_j_15;	// matmul/matmul-hw.mlir:23252:23
  wire [31:0]     b_i_k_6_i_j_15;	// matmul/matmul-hw.mlir:23255:23
  wire [31:0]     c_prev_i_k_6_i_j_15;	// matmul/matmul-hw.mlir:23258:28
  wire            tk_i_k_6_i_j_15;	// matmul/matmul-hw.mlir:23261:24
  wire [31:0]     c_i_k_6_i_j_15;	// matmul/matmul-hw.mlir:23265:23
  reg  [3:0]      i_k_next_4028;	// matmul/matmul-hw.mlir:23270:22
  wire [31:0]     a_i_k_7_i_j_15;	// matmul/matmul-hw.mlir:23282:23
  wire [31:0]     b_i_k_7_i_j_15;	// matmul/matmul-hw.mlir:23285:23
  wire [31:0]     c_prev_i_k_7_i_j_15;	// matmul/matmul-hw.mlir:23288:28
  wire            tk_i_k_7_i_j_15;	// matmul/matmul-hw.mlir:23291:24
  wire [31:0]     c_i_k_7_i_j_15;	// matmul/matmul-hw.mlir:23295:23
  reg  [3:0]      i_k_next_4031;	// matmul/matmul-hw.mlir:23300:22
  wire [31:0]     a_i_k_8_i_j_15;	// matmul/matmul-hw.mlir:23312:23
  wire [31:0]     b_i_k_8_i_j_15;	// matmul/matmul-hw.mlir:23315:23
  wire [31:0]     c_prev_i_k_8_i_j_15;	// matmul/matmul-hw.mlir:23318:28
  wire            tk_i_k_8_i_j_15;	// matmul/matmul-hw.mlir:23321:24
  wire [31:0]     c_i_k_8_i_j_15;	// matmul/matmul-hw.mlir:23325:23
  reg  [3:0]      i_k_next_4034;	// matmul/matmul-hw.mlir:23330:22
  wire [31:0]     a_i_k_9_i_j_15;	// matmul/matmul-hw.mlir:23342:23
  wire [31:0]     b_i_k_9_i_j_15;	// matmul/matmul-hw.mlir:23345:23
  wire [31:0]     c_prev_i_k_9_i_j_15;	// matmul/matmul-hw.mlir:23348:28
  wire            tk_i_k_9_i_j_15;	// matmul/matmul-hw.mlir:23351:24
  wire [31:0]     c_i_k_9_i_j_15;	// matmul/matmul-hw.mlir:23355:23
  reg  [3:0]      i_k_next_4037;	// matmul/matmul-hw.mlir:23360:22
  wire [31:0]     a_i_k_10_i_j_15;	// matmul/matmul-hw.mlir:23372:24
  wire [31:0]     b_i_k_10_i_j_15;	// matmul/matmul-hw.mlir:23375:24
  wire [31:0]     c_prev_i_k_10_i_j_15;	// matmul/matmul-hw.mlir:23378:29
  wire            tk_i_k_10_i_j_15;	// matmul/matmul-hw.mlir:23381:25
  wire [31:0]     c_i_k_10_i_j_15;	// matmul/matmul-hw.mlir:23385:24
  reg  [3:0]      i_k_next_4040;	// matmul/matmul-hw.mlir:23390:22
  wire [31:0]     a_i_k_11_i_j_15;	// matmul/matmul-hw.mlir:23402:24
  wire [31:0]     b_i_k_11_i_j_15;	// matmul/matmul-hw.mlir:23405:24
  wire [31:0]     c_prev_i_k_11_i_j_15;	// matmul/matmul-hw.mlir:23408:29
  wire            tk_i_k_11_i_j_15;	// matmul/matmul-hw.mlir:23411:25
  wire [31:0]     c_i_k_11_i_j_15;	// matmul/matmul-hw.mlir:23415:24
  reg  [3:0]      i_k_next_4043;	// matmul/matmul-hw.mlir:23420:22
  wire [31:0]     a_i_k_12_i_j_15;	// matmul/matmul-hw.mlir:23432:24
  wire [31:0]     b_i_k_12_i_j_15;	// matmul/matmul-hw.mlir:23435:24
  wire [31:0]     c_prev_i_k_12_i_j_15;	// matmul/matmul-hw.mlir:23438:29
  wire            tk_i_k_12_i_j_15;	// matmul/matmul-hw.mlir:23441:25
  wire [31:0]     c_i_k_12_i_j_15;	// matmul/matmul-hw.mlir:23445:24
  reg  [3:0]      i_k_next_4046;	// matmul/matmul-hw.mlir:23450:22
  wire [31:0]     a_i_k_13_i_j_15;	// matmul/matmul-hw.mlir:23462:24
  wire [31:0]     b_i_k_13_i_j_15;	// matmul/matmul-hw.mlir:23465:24
  wire [31:0]     c_prev_i_k_13_i_j_15;	// matmul/matmul-hw.mlir:23468:29
  wire            tk_i_k_13_i_j_15;	// matmul/matmul-hw.mlir:23471:25
  wire [31:0]     c_i_k_13_i_j_15;	// matmul/matmul-hw.mlir:23475:24
  reg  [3:0]      i_k_next_4049;	// matmul/matmul-hw.mlir:23480:22
  wire [31:0]     a_i_k_14_i_j_15;	// matmul/matmul-hw.mlir:23492:24
  wire [31:0]     b_i_k_14_i_j_15;	// matmul/matmul-hw.mlir:23495:24
  wire [31:0]     c_prev_i_k_14_i_j_15;	// matmul/matmul-hw.mlir:23498:29
  wire            tk_i_k_14_i_j_15;	// matmul/matmul-hw.mlir:23501:25
  wire [31:0]     c_i_k_14_i_j_15;	// matmul/matmul-hw.mlir:23505:24
  reg  [3:0]      i_k_next_4052;	// matmul/matmul-hw.mlir:23510:22
  wire [31:0]     a_i_k_15_i_j_15;	// matmul/matmul-hw.mlir:23522:24
  wire [31:0]     b_i_k_15_i_j_15;	// matmul/matmul-hw.mlir:23525:24
  wire [31:0]     c_prev_i_k_15_i_j_15;	// matmul/matmul-hw.mlir:23528:29
  wire            tk_i_k_15_i_j_15;	// matmul/matmul-hw.mlir:23531:25
  wire [31:0]     c_i_k_15_i_j_15;	// matmul/matmul-hw.mlir:23535:24
  reg  [3:0]      i_k_next_4055;	// matmul/matmul-hw.mlir:23540:22
  reg  [34:0]     _T_4057;	// matmul/matmul-hw.mlir:23548:13
  reg  [3:0][3:0] i_delayed_4062;	// matmul/matmul-hw.mlir:23564:23

  wire [31:0] _T_2454 = B_p0_rd_data[8'h0];	// matmul/matmul-hw.mlir:10297:14, :10298:10
  wire [31:0] _T_2455 = B_p0_rd_data[8'h1];	// matmul/matmul-hw.mlir:10300:14, :10301:10
  wire [31:0] _T_2456 = B_p0_rd_data[8'h2];	// matmul/matmul-hw.mlir:10303:14, :10304:11
  wire [31:0] _T_2457 = B_p0_rd_data[8'h3];	// matmul/matmul-hw.mlir:10306:14, :10307:11
  wire [31:0] _T_2458 = B_p0_rd_data[8'h4];	// matmul/matmul-hw.mlir:10309:14, :10310:11
  wire [31:0] _T_2459 = B_p0_rd_data[8'h5];	// matmul/matmul-hw.mlir:10312:14, :10313:11
  wire [31:0] _T_2460 = B_p0_rd_data[8'h6];	// matmul/matmul-hw.mlir:10315:14, :10316:11
  wire [31:0] _T_2461 = B_p0_rd_data[8'h7];	// matmul/matmul-hw.mlir:10318:14, :10319:11
  wire [31:0] _T_2462 = B_p0_rd_data[8'h8];	// matmul/matmul-hw.mlir:10321:14, :10322:11
  wire [31:0] _T_2463 = B_p0_rd_data[8'h9];	// matmul/matmul-hw.mlir:10324:14, :10325:11
  wire [31:0] _T_2464 = B_p0_rd_data[8'hA];	// matmul/matmul-hw.mlir:10327:15, :10328:11
  wire [31:0] _T_2465 = B_p0_rd_data[8'hB];	// matmul/matmul-hw.mlir:10330:15, :10331:11
  wire [31:0] _T_2466 = B_p0_rd_data[8'hC];	// matmul/matmul-hw.mlir:10333:15, :10334:11
  wire [31:0] _T_2467 = B_p0_rd_data[8'hD];	// matmul/matmul-hw.mlir:10336:15, :10337:11
  wire [31:0] _T_2468 = B_p0_rd_data[8'hE];	// matmul/matmul-hw.mlir:10339:15, :10340:11
  wire [31:0] _T_2469 = B_p0_rd_data[8'hF];	// matmul/matmul-hw.mlir:10342:15, :10343:11
  wire [31:0] _T_2470 = B_p0_rd_data[8'h10];	// matmul/matmul-hw.mlir:10345:15, :10346:11
  wire [31:0] _T_2471 = B_p0_rd_data[8'h11];	// matmul/matmul-hw.mlir:10348:15, :10349:11
  wire [31:0] _T_2472 = B_p0_rd_data[8'h12];	// matmul/matmul-hw.mlir:10351:15, :10352:11
  wire [31:0] _T_2473 = B_p0_rd_data[8'h13];	// matmul/matmul-hw.mlir:10354:15, :10355:11
  wire [31:0] _T_2474 = B_p0_rd_data[8'h14];	// matmul/matmul-hw.mlir:10357:15, :10358:11
  wire [31:0] _T_2475 = B_p0_rd_data[8'h15];	// matmul/matmul-hw.mlir:10360:15, :10361:11
  wire [31:0] _T_2476 = B_p0_rd_data[8'h16];	// matmul/matmul-hw.mlir:10363:15, :10364:11
  wire [31:0] _T_2477 = B_p0_rd_data[8'h17];	// matmul/matmul-hw.mlir:10366:15, :10367:11
  wire [31:0] _T_2478 = B_p0_rd_data[8'h18];	// matmul/matmul-hw.mlir:10369:15, :10370:11
  wire [31:0] _T_2479 = B_p0_rd_data[8'h19];	// matmul/matmul-hw.mlir:10372:15, :10373:11
  wire [31:0] _T_2480 = B_p0_rd_data[8'h1A];	// matmul/matmul-hw.mlir:10375:15, :10376:11
  wire [31:0] _T_2481 = B_p0_rd_data[8'h1B];	// matmul/matmul-hw.mlir:10378:15, :10379:11
  wire [31:0] _T_2482 = B_p0_rd_data[8'h1C];	// matmul/matmul-hw.mlir:10381:15, :10382:11
  wire [31:0] _T_2483 = B_p0_rd_data[8'h1D];	// matmul/matmul-hw.mlir:10384:15, :10385:11
  wire [31:0] _T_2484 = B_p0_rd_data[8'h1E];	// matmul/matmul-hw.mlir:10387:15, :10388:11
  wire [31:0] _T_2485 = B_p0_rd_data[8'h1F];	// matmul/matmul-hw.mlir:10390:15, :10391:11
  wire [31:0] _T_2486 = B_p0_rd_data[8'h20];	// matmul/matmul-hw.mlir:10393:15, :10394:11
  wire [31:0] _T_2487 = B_p0_rd_data[8'h21];	// matmul/matmul-hw.mlir:10396:15, :10397:11
  wire [31:0] _T_2488 = B_p0_rd_data[8'h22];	// matmul/matmul-hw.mlir:10399:15, :10400:11
  wire [31:0] _T_2489 = B_p0_rd_data[8'h23];	// matmul/matmul-hw.mlir:10402:15, :10403:11
  wire [31:0] _T_2490 = B_p0_rd_data[8'h24];	// matmul/matmul-hw.mlir:10405:15, :10406:11
  wire [31:0] _T_2491 = B_p0_rd_data[8'h25];	// matmul/matmul-hw.mlir:10408:15, :10409:11
  wire [31:0] _T_2492 = B_p0_rd_data[8'h26];	// matmul/matmul-hw.mlir:10411:15, :10412:11
  wire [31:0] _T_2493 = B_p0_rd_data[8'h27];	// matmul/matmul-hw.mlir:10414:15, :10415:11
  wire [31:0] _T_2494 = B_p0_rd_data[8'h28];	// matmul/matmul-hw.mlir:10417:15, :10418:11
  wire [31:0] _T_2495 = B_p0_rd_data[8'h29];	// matmul/matmul-hw.mlir:10420:15, :10421:11
  wire [31:0] _T_2496 = B_p0_rd_data[8'h2A];	// matmul/matmul-hw.mlir:10423:15, :10424:11
  wire [31:0] _T_2497 = B_p0_rd_data[8'h2B];	// matmul/matmul-hw.mlir:10426:15, :10427:11
  wire [31:0] _T_2498 = B_p0_rd_data[8'h2C];	// matmul/matmul-hw.mlir:10429:15, :10430:11
  wire [31:0] _T_2499 = B_p0_rd_data[8'h2D];	// matmul/matmul-hw.mlir:10432:15, :10433:11
  wire [31:0] _T_2500 = B_p0_rd_data[8'h2E];	// matmul/matmul-hw.mlir:10435:15, :10436:11
  wire [31:0] _T_2501 = B_p0_rd_data[8'h2F];	// matmul/matmul-hw.mlir:10438:15, :10439:11
  wire [31:0] _T_2502 = B_p0_rd_data[8'h30];	// matmul/matmul-hw.mlir:10441:15, :10442:11
  wire [31:0] _T_2503 = B_p0_rd_data[8'h31];	// matmul/matmul-hw.mlir:10444:15, :10445:11
  wire [31:0] _T_2504 = B_p0_rd_data[8'h32];	// matmul/matmul-hw.mlir:10447:15, :10448:11
  wire [31:0] _T_2505 = B_p0_rd_data[8'h33];	// matmul/matmul-hw.mlir:10450:15, :10451:11
  wire [31:0] _T_2506 = B_p0_rd_data[8'h34];	// matmul/matmul-hw.mlir:10453:15, :10454:11
  wire [31:0] _T_2507 = B_p0_rd_data[8'h35];	// matmul/matmul-hw.mlir:10456:15, :10457:11
  wire [31:0] _T_2508 = B_p0_rd_data[8'h36];	// matmul/matmul-hw.mlir:10459:15, :10460:11
  wire [31:0] _T_2509 = B_p0_rd_data[8'h37];	// matmul/matmul-hw.mlir:10462:15, :10463:11
  wire [31:0] _T_2510 = B_p0_rd_data[8'h38];	// matmul/matmul-hw.mlir:10465:15, :10466:11
  wire [31:0] _T_2511 = B_p0_rd_data[8'h39];	// matmul/matmul-hw.mlir:10468:15, :10469:11
  wire [31:0] _T_2512 = B_p0_rd_data[8'h3A];	// matmul/matmul-hw.mlir:10471:15, :10472:11
  wire [31:0] _T_2513 = B_p0_rd_data[8'h3B];	// matmul/matmul-hw.mlir:10474:15, :10475:11
  wire [31:0] _T_2514 = B_p0_rd_data[8'h3C];	// matmul/matmul-hw.mlir:10477:15, :10478:11
  wire [31:0] _T_2515 = B_p0_rd_data[8'h3D];	// matmul/matmul-hw.mlir:10480:15, :10481:11
  wire [31:0] _T_2516 = B_p0_rd_data[8'h3E];	// matmul/matmul-hw.mlir:10483:15, :10484:11
  wire [31:0] _T_2517 = B_p0_rd_data[8'h3F];	// matmul/matmul-hw.mlir:10486:15, :10487:11
  wire [31:0] _T_2518 = B_p0_rd_data[8'h40];	// matmul/matmul-hw.mlir:10489:15, :10490:11
  wire [31:0] _T_2519 = B_p0_rd_data[8'h41];	// matmul/matmul-hw.mlir:10492:15, :10493:11
  wire [31:0] _T_2520 = B_p0_rd_data[8'h42];	// matmul/matmul-hw.mlir:10495:15, :10496:11
  wire [31:0] _T_2521 = B_p0_rd_data[8'h43];	// matmul/matmul-hw.mlir:10498:15, :10499:11
  wire [31:0] _T_2522 = B_p0_rd_data[8'h44];	// matmul/matmul-hw.mlir:10501:15, :10502:11
  wire [31:0] _T_2523 = B_p0_rd_data[8'h45];	// matmul/matmul-hw.mlir:10504:15, :10505:11
  wire [31:0] _T_2524 = B_p0_rd_data[8'h46];	// matmul/matmul-hw.mlir:10507:15, :10508:11
  wire [31:0] _T_2525 = B_p0_rd_data[8'h47];	// matmul/matmul-hw.mlir:10510:15, :10511:11
  wire [31:0] _T_2526 = B_p0_rd_data[8'h48];	// matmul/matmul-hw.mlir:10513:15, :10514:11
  wire [31:0] _T_2527 = B_p0_rd_data[8'h49];	// matmul/matmul-hw.mlir:10516:15, :10517:11
  wire [31:0] _T_2528 = B_p0_rd_data[8'h4A];	// matmul/matmul-hw.mlir:10519:15, :10520:11
  wire [31:0] _T_2529 = B_p0_rd_data[8'h4B];	// matmul/matmul-hw.mlir:10522:15, :10523:11
  wire [31:0] _T_2530 = B_p0_rd_data[8'h4C];	// matmul/matmul-hw.mlir:10525:15, :10526:11
  wire [31:0] _T_2531 = B_p0_rd_data[8'h4D];	// matmul/matmul-hw.mlir:10528:15, :10529:11
  wire [31:0] _T_2532 = B_p0_rd_data[8'h4E];	// matmul/matmul-hw.mlir:10531:15, :10532:11
  wire [31:0] _T_2533 = B_p0_rd_data[8'h4F];	// matmul/matmul-hw.mlir:10534:15, :10535:11
  wire [31:0] _T_2534 = B_p0_rd_data[8'h50];	// matmul/matmul-hw.mlir:10537:15, :10538:11
  wire [31:0] _T_2535 = B_p0_rd_data[8'h51];	// matmul/matmul-hw.mlir:10540:15, :10541:11
  wire [31:0] _T_2536 = B_p0_rd_data[8'h52];	// matmul/matmul-hw.mlir:10543:15, :10544:11
  wire [31:0] _T_2537 = B_p0_rd_data[8'h53];	// matmul/matmul-hw.mlir:10546:15, :10547:11
  wire [31:0] _T_2538 = B_p0_rd_data[8'h54];	// matmul/matmul-hw.mlir:10549:15, :10550:11
  wire [31:0] _T_2539 = B_p0_rd_data[8'h55];	// matmul/matmul-hw.mlir:10552:15, :10553:11
  wire [31:0] _T_2540 = B_p0_rd_data[8'h56];	// matmul/matmul-hw.mlir:10555:15, :10556:11
  wire [31:0] _T_2541 = B_p0_rd_data[8'h57];	// matmul/matmul-hw.mlir:10558:15, :10559:11
  wire [31:0] _T_2542 = B_p0_rd_data[8'h58];	// matmul/matmul-hw.mlir:10561:15, :10562:11
  wire [31:0] _T_2543 = B_p0_rd_data[8'h59];	// matmul/matmul-hw.mlir:10564:15, :10565:11
  wire [31:0] _T_2544 = B_p0_rd_data[8'h5A];	// matmul/matmul-hw.mlir:10567:15, :10568:11
  wire [31:0] _T_2545 = B_p0_rd_data[8'h5B];	// matmul/matmul-hw.mlir:10570:15, :10571:11
  wire [31:0] _T_2546 = B_p0_rd_data[8'h5C];	// matmul/matmul-hw.mlir:10573:15, :10574:12
  wire [31:0] _T_2547 = B_p0_rd_data[8'h5D];	// matmul/matmul-hw.mlir:10576:15, :10577:12
  wire [31:0] _T_2548 = B_p0_rd_data[8'h5E];	// matmul/matmul-hw.mlir:10579:15, :10580:12
  wire [31:0] _T_2549 = B_p0_rd_data[8'h5F];	// matmul/matmul-hw.mlir:10582:15, :10583:12
  wire [31:0] _T_2550 = B_p0_rd_data[8'h60];	// matmul/matmul-hw.mlir:10585:15, :10586:12
  wire [31:0] _T_2551 = B_p0_rd_data[8'h61];	// matmul/matmul-hw.mlir:10588:15, :10589:12
  wire [31:0] _T_2552 = B_p0_rd_data[8'h62];	// matmul/matmul-hw.mlir:10591:15, :10592:12
  wire [31:0] _T_2553 = B_p0_rd_data[8'h63];	// matmul/matmul-hw.mlir:10594:15, :10595:12
  wire [31:0] _T_2554 = B_p0_rd_data[8'h64];	// matmul/matmul-hw.mlir:10597:16, :10598:12
  wire [31:0] _T_2555 = B_p0_rd_data[8'h65];	// matmul/matmul-hw.mlir:10600:16, :10601:12
  wire [31:0] _T_2556 = B_p0_rd_data[8'h66];	// matmul/matmul-hw.mlir:10603:16, :10604:12
  wire [31:0] _T_2557 = B_p0_rd_data[8'h67];	// matmul/matmul-hw.mlir:10606:16, :10607:12
  wire [31:0] _T_2558 = B_p0_rd_data[8'h68];	// matmul/matmul-hw.mlir:10609:16, :10610:12
  wire [31:0] _T_2559 = B_p0_rd_data[8'h69];	// matmul/matmul-hw.mlir:10612:16, :10613:12
  wire [31:0] _T_2560 = B_p0_rd_data[8'h6A];	// matmul/matmul-hw.mlir:10615:16, :10616:12
  wire [31:0] _T_2561 = B_p0_rd_data[8'h6B];	// matmul/matmul-hw.mlir:10618:16, :10619:12
  wire [31:0] _T_2562 = B_p0_rd_data[8'h6C];	// matmul/matmul-hw.mlir:10621:16, :10622:12
  wire [31:0] _T_2563 = B_p0_rd_data[8'h6D];	// matmul/matmul-hw.mlir:10624:16, :10625:12
  wire [31:0] _T_2564 = B_p0_rd_data[8'h6E];	// matmul/matmul-hw.mlir:10627:16, :10628:12
  wire [31:0] _T_2565 = B_p0_rd_data[8'h6F];	// matmul/matmul-hw.mlir:10630:16, :10631:12
  wire [31:0] _T_2566 = B_p0_rd_data[8'h70];	// matmul/matmul-hw.mlir:10633:16, :10634:12
  wire [31:0] _T_2567 = B_p0_rd_data[8'h71];	// matmul/matmul-hw.mlir:10636:16, :10637:12
  wire [31:0] _T_2568 = B_p0_rd_data[8'h72];	// matmul/matmul-hw.mlir:10639:16, :10640:12
  wire [31:0] _T_2569 = B_p0_rd_data[8'h73];	// matmul/matmul-hw.mlir:10642:16, :10643:12
  wire [31:0] _T_2570 = B_p0_rd_data[8'h74];	// matmul/matmul-hw.mlir:10645:16, :10646:12
  wire [31:0] _T_2571 = B_p0_rd_data[8'h75];	// matmul/matmul-hw.mlir:10648:16, :10649:12
  wire [31:0] _T_2572 = B_p0_rd_data[8'h76];	// matmul/matmul-hw.mlir:10651:16, :10652:12
  wire [31:0] _T_2573 = B_p0_rd_data[8'h77];	// matmul/matmul-hw.mlir:10654:16, :10655:12
  wire [31:0] _T_2574 = B_p0_rd_data[8'h78];	// matmul/matmul-hw.mlir:10657:16, :10658:12
  wire [31:0] _T_2575 = B_p0_rd_data[8'h79];	// matmul/matmul-hw.mlir:10660:16, :10661:12
  wire [31:0] _T_2576 = B_p0_rd_data[8'h7A];	// matmul/matmul-hw.mlir:10663:16, :10664:12
  wire [31:0] _T_2577 = B_p0_rd_data[8'h7B];	// matmul/matmul-hw.mlir:10666:16, :10667:12
  wire [31:0] _T_2578 = B_p0_rd_data[8'h7C];	// matmul/matmul-hw.mlir:10669:16, :10670:12
  wire [31:0] _T_2579 = B_p0_rd_data[8'h7D];	// matmul/matmul-hw.mlir:10672:16, :10673:12
  wire [31:0] _T_2580 = B_p0_rd_data[8'h7E];	// matmul/matmul-hw.mlir:10675:16, :10676:12
  wire [31:0] _T_2581 = B_p0_rd_data[8'h7F];	// matmul/matmul-hw.mlir:10678:16, :10679:12
  wire [31:0] _T_2582 = B_p0_rd_data[8'h80];	// matmul/matmul-hw.mlir:10681:17, :10682:12
  wire [31:0] _T_2583 = B_p0_rd_data[8'h81];	// matmul/matmul-hw.mlir:10684:17, :10685:12
  wire [31:0] _T_2584 = B_p0_rd_data[8'h82];	// matmul/matmul-hw.mlir:10687:17, :10688:12
  wire [31:0] _T_2585 = B_p0_rd_data[8'h83];	// matmul/matmul-hw.mlir:10690:17, :10691:12
  wire [31:0] _T_2586 = B_p0_rd_data[8'h84];	// matmul/matmul-hw.mlir:10693:17, :10694:12
  wire [31:0] _T_2587 = B_p0_rd_data[8'h85];	// matmul/matmul-hw.mlir:10696:17, :10697:12
  wire [31:0] _T_2588 = B_p0_rd_data[8'h86];	// matmul/matmul-hw.mlir:10699:17, :10700:12
  wire [31:0] _T_2589 = B_p0_rd_data[8'h87];	// matmul/matmul-hw.mlir:10702:17, :10703:12
  wire [31:0] _T_2590 = B_p0_rd_data[8'h88];	// matmul/matmul-hw.mlir:10705:17, :10706:12
  wire [31:0] _T_2591 = B_p0_rd_data[8'h89];	// matmul/matmul-hw.mlir:10708:17, :10709:12
  wire [31:0] _T_2592 = B_p0_rd_data[8'h8A];	// matmul/matmul-hw.mlir:10711:17, :10712:12
  wire [31:0] _T_2593 = B_p0_rd_data[8'h8B];	// matmul/matmul-hw.mlir:10714:17, :10715:12
  wire [31:0] _T_2594 = B_p0_rd_data[8'h8C];	// matmul/matmul-hw.mlir:10717:17, :10718:12
  wire [31:0] _T_2595 = B_p0_rd_data[8'h8D];	// matmul/matmul-hw.mlir:10720:17, :10721:12
  wire [31:0] _T_2596 = B_p0_rd_data[8'h8E];	// matmul/matmul-hw.mlir:10723:17, :10724:12
  wire [31:0] _T_2597 = B_p0_rd_data[8'h8F];	// matmul/matmul-hw.mlir:10726:17, :10727:12
  wire [31:0] _T_2598 = B_p0_rd_data[8'h90];	// matmul/matmul-hw.mlir:10729:17, :10730:12
  wire [31:0] _T_2599 = B_p0_rd_data[8'h91];	// matmul/matmul-hw.mlir:10732:17, :10733:12
  wire [31:0] _T_2600 = B_p0_rd_data[8'h92];	// matmul/matmul-hw.mlir:10735:17, :10736:12
  wire [31:0] _T_2601 = B_p0_rd_data[8'h93];	// matmul/matmul-hw.mlir:10738:17, :10739:12
  wire [31:0] _T_2602 = B_p0_rd_data[8'h94];	// matmul/matmul-hw.mlir:10741:17, :10742:12
  wire [31:0] _T_2603 = B_p0_rd_data[8'h95];	// matmul/matmul-hw.mlir:10744:17, :10745:12
  wire [31:0] _T_2604 = B_p0_rd_data[8'h96];	// matmul/matmul-hw.mlir:10747:17, :10748:12
  wire [31:0] _T_2605 = B_p0_rd_data[8'h97];	// matmul/matmul-hw.mlir:10750:17, :10751:12
  wire [31:0] _T_2606 = B_p0_rd_data[8'h98];	// matmul/matmul-hw.mlir:10753:17, :10754:12
  wire [31:0] _T_2607 = B_p0_rd_data[8'h99];	// matmul/matmul-hw.mlir:10756:17, :10757:12
  wire [31:0] _T_2608 = B_p0_rd_data[8'h9A];	// matmul/matmul-hw.mlir:10759:17, :10760:12
  wire [31:0] _T_2609 = B_p0_rd_data[8'h9B];	// matmul/matmul-hw.mlir:10762:17, :10763:12
  wire [31:0] _T_2610 = B_p0_rd_data[8'h9C];	// matmul/matmul-hw.mlir:10765:17, :10766:12
  wire [31:0] _T_2611 = B_p0_rd_data[8'h9D];	// matmul/matmul-hw.mlir:10768:16, :10769:12
  wire [31:0] _T_2612 = B_p0_rd_data[8'h9E];	// matmul/matmul-hw.mlir:10771:16, :10772:12
  wire [31:0] _T_2613 = B_p0_rd_data[8'h9F];	// matmul/matmul-hw.mlir:10774:16, :10775:12
  wire [31:0] _T_2614 = B_p0_rd_data[8'hA0];	// matmul/matmul-hw.mlir:10777:16, :10778:12
  wire [31:0] _T_2615 = B_p0_rd_data[8'hA1];	// matmul/matmul-hw.mlir:10780:16, :10781:12
  wire [31:0] _T_2616 = B_p0_rd_data[8'hA2];	// matmul/matmul-hw.mlir:10783:16, :10784:12
  wire [31:0] _T_2617 = B_p0_rd_data[8'hA3];	// matmul/matmul-hw.mlir:10786:16, :10787:12
  wire [31:0] _T_2618 = B_p0_rd_data[8'hA4];	// matmul/matmul-hw.mlir:10789:16, :10790:12
  wire [31:0] _T_2619 = B_p0_rd_data[8'hA5];	// matmul/matmul-hw.mlir:10792:16, :10793:12
  wire [31:0] _T_2620 = B_p0_rd_data[8'hA6];	// matmul/matmul-hw.mlir:10795:16, :10796:12
  wire [31:0] _T_2621 = B_p0_rd_data[8'hA7];	// matmul/matmul-hw.mlir:10798:16, :10799:12
  wire [31:0] _T_2622 = B_p0_rd_data[8'hA8];	// matmul/matmul-hw.mlir:10801:16, :10802:12
  wire [31:0] _T_2623 = B_p0_rd_data[8'hA9];	// matmul/matmul-hw.mlir:10804:16, :10805:12
  wire [31:0] _T_2624 = B_p0_rd_data[8'hAA];	// matmul/matmul-hw.mlir:10807:16, :10808:12
  wire [31:0] _T_2625 = B_p0_rd_data[8'hAB];	// matmul/matmul-hw.mlir:10810:16, :10811:12
  wire [31:0] _T_2626 = B_p0_rd_data[8'hAC];	// matmul/matmul-hw.mlir:10813:16, :10814:12
  wire [31:0] _T_2627 = B_p0_rd_data[8'hAD];	// matmul/matmul-hw.mlir:10816:16, :10817:12
  wire [31:0] _T_2628 = B_p0_rd_data[8'hAE];	// matmul/matmul-hw.mlir:10819:16, :10820:12
  wire [31:0] _T_2629 = B_p0_rd_data[8'hAF];	// matmul/matmul-hw.mlir:10822:16, :10823:12
  wire [31:0] _T_2630 = B_p0_rd_data[8'hB0];	// matmul/matmul-hw.mlir:10825:16, :10826:12
  wire [31:0] _T_2631 = B_p0_rd_data[8'hB1];	// matmul/matmul-hw.mlir:10828:16, :10829:12
  wire [31:0] _T_2632 = B_p0_rd_data[8'hB2];	// matmul/matmul-hw.mlir:10831:16, :10832:12
  wire [31:0] _T_2633 = B_p0_rd_data[8'hB3];	// matmul/matmul-hw.mlir:10834:16, :10835:12
  wire [31:0] _T_2634 = B_p0_rd_data[8'hB4];	// matmul/matmul-hw.mlir:10837:16, :10838:12
  wire [31:0] _T_2635 = B_p0_rd_data[8'hB5];	// matmul/matmul-hw.mlir:10840:16, :10841:12
  wire [31:0] _T_2636 = B_p0_rd_data[8'hB6];	// matmul/matmul-hw.mlir:10843:16, :10844:12
  wire [31:0] _T_2637 = B_p0_rd_data[8'hB7];	// matmul/matmul-hw.mlir:10846:16, :10847:12
  wire [31:0] _T_2638 = B_p0_rd_data[8'hB8];	// matmul/matmul-hw.mlir:10849:16, :10850:12
  wire [31:0] _T_2639 = B_p0_rd_data[8'hB9];	// matmul/matmul-hw.mlir:10852:16, :10853:12
  wire [31:0] _T_2640 = B_p0_rd_data[8'hBA];	// matmul/matmul-hw.mlir:10855:16, :10856:12
  wire [31:0] _T_2641 = B_p0_rd_data[8'hBB];	// matmul/matmul-hw.mlir:10858:16, :10859:12
  wire [31:0] _T_2642 = B_p0_rd_data[8'hBC];	// matmul/matmul-hw.mlir:10861:16, :10862:12
  wire [31:0] _T_2643 = B_p0_rd_data[8'hBD];	// matmul/matmul-hw.mlir:10864:16, :10865:12
  wire [31:0] _T_2644 = B_p0_rd_data[8'hBE];	// matmul/matmul-hw.mlir:10867:16, :10868:12
  wire [31:0] _T_2645 = B_p0_rd_data[8'hBF];	// matmul/matmul-hw.mlir:10870:16, :10871:12
  wire [31:0] _T_2646 = B_p0_rd_data[8'hC0];	// matmul/matmul-hw.mlir:10873:16, :10874:12
  wire [31:0] _T_2647 = B_p0_rd_data[8'hC1];	// matmul/matmul-hw.mlir:10876:16, :10877:12
  wire [31:0] _T_2648 = B_p0_rd_data[8'hC2];	// matmul/matmul-hw.mlir:10879:16, :10880:12
  wire [31:0] _T_2649 = B_p0_rd_data[8'hC3];	// matmul/matmul-hw.mlir:10882:16, :10883:12
  wire [31:0] _T_2650 = B_p0_rd_data[8'hC4];	// matmul/matmul-hw.mlir:10885:16, :10886:12
  wire [31:0] _T_2651 = B_p0_rd_data[8'hC5];	// matmul/matmul-hw.mlir:10888:16, :10889:12
  wire [31:0] _T_2652 = B_p0_rd_data[8'hC6];	// matmul/matmul-hw.mlir:10891:16, :10892:12
  wire [31:0] _T_2653 = B_p0_rd_data[8'hC7];	// matmul/matmul-hw.mlir:10894:16, :10895:12
  wire [31:0] _T_2654 = B_p0_rd_data[8'hC8];	// matmul/matmul-hw.mlir:10897:16, :10898:12
  wire [31:0] _T_2655 = B_p0_rd_data[8'hC9];	// matmul/matmul-hw.mlir:10900:16, :10901:12
  wire [31:0] _T_2656 = B_p0_rd_data[8'hCA];	// matmul/matmul-hw.mlir:10903:16, :10904:12
  wire [31:0] _T_2657 = B_p0_rd_data[8'hCB];	// matmul/matmul-hw.mlir:10906:16, :10907:12
  wire [31:0] _T_2658 = B_p0_rd_data[8'hCC];	// matmul/matmul-hw.mlir:10909:16, :10910:12
  wire [31:0] _T_2659 = B_p0_rd_data[8'hCD];	// matmul/matmul-hw.mlir:10912:16, :10913:12
  wire [31:0] _T_2660 = B_p0_rd_data[8'hCE];	// matmul/matmul-hw.mlir:10915:16, :10916:12
  wire [31:0] _T_2661 = B_p0_rd_data[8'hCF];	// matmul/matmul-hw.mlir:10918:16, :10919:12
  wire [31:0] _T_2662 = B_p0_rd_data[8'hD0];	// matmul/matmul-hw.mlir:10921:16, :10922:12
  wire [31:0] _T_2663 = B_p0_rd_data[8'hD1];	// matmul/matmul-hw.mlir:10924:16, :10925:12
  wire [31:0] _T_2664 = B_p0_rd_data[8'hD2];	// matmul/matmul-hw.mlir:10927:16, :10928:12
  wire [31:0] _T_2665 = B_p0_rd_data[8'hD3];	// matmul/matmul-hw.mlir:10930:16, :10931:12
  wire [31:0] _T_2666 = B_p0_rd_data[8'hD4];	// matmul/matmul-hw.mlir:10933:16, :10934:12
  wire [31:0] _T_2667 = B_p0_rd_data[8'hD5];	// matmul/matmul-hw.mlir:10936:16, :10937:12
  wire [31:0] _T_2668 = B_p0_rd_data[8'hD6];	// matmul/matmul-hw.mlir:10939:16, :10940:12
  wire [31:0] _T_2669 = B_p0_rd_data[8'hD7];	// matmul/matmul-hw.mlir:10942:16, :10943:12
  wire [31:0] _T_2670 = B_p0_rd_data[8'hD8];	// matmul/matmul-hw.mlir:10945:16, :10946:12
  wire [31:0] _T_2671 = B_p0_rd_data[8'hD9];	// matmul/matmul-hw.mlir:10948:16, :10949:12
  wire [31:0] _T_2672 = B_p0_rd_data[8'hDA];	// matmul/matmul-hw.mlir:10951:16, :10952:12
  wire [31:0] _T_2673 = B_p0_rd_data[8'hDB];	// matmul/matmul-hw.mlir:10954:16, :10955:12
  wire [31:0] _T_2674 = B_p0_rd_data[8'hDC];	// matmul/matmul-hw.mlir:10957:16, :10958:12
  wire [31:0] _T_2675 = B_p0_rd_data[8'hDD];	// matmul/matmul-hw.mlir:10960:16, :10961:12
  wire [31:0] _T_2676 = B_p0_rd_data[8'hDE];	// matmul/matmul-hw.mlir:10963:16, :10964:12
  wire [31:0] _T_2677 = B_p0_rd_data[8'hDF];	// matmul/matmul-hw.mlir:10966:16, :10967:12
  wire [31:0] _T_2678 = B_p0_rd_data[8'hE0];	// matmul/matmul-hw.mlir:10969:16, :10970:12
  wire [31:0] _T_2679 = B_p0_rd_data[8'hE1];	// matmul/matmul-hw.mlir:10972:16, :10973:12
  wire [31:0] _T_2680 = B_p0_rd_data[8'hE2];	// matmul/matmul-hw.mlir:10975:16, :10976:12
  wire [31:0] _T_2681 = B_p0_rd_data[8'hE3];	// matmul/matmul-hw.mlir:10978:16, :10979:12
  wire [31:0] _T_2682 = B_p0_rd_data[8'hE4];	// matmul/matmul-hw.mlir:10981:16, :10982:12
  wire [31:0] _T_2683 = B_p0_rd_data[8'hE5];	// matmul/matmul-hw.mlir:10984:16, :10985:12
  wire [31:0] _T_2684 = B_p0_rd_data[8'hE6];	// matmul/matmul-hw.mlir:10987:16, :10988:12
  wire [31:0] _T_2685 = B_p0_rd_data[8'hE7];	// matmul/matmul-hw.mlir:10990:16, :10991:12
  wire [31:0] _T_2686 = B_p0_rd_data[8'hE8];	// matmul/matmul-hw.mlir:10993:16, :10994:12
  wire [31:0] _T_2687 = B_p0_rd_data[8'hE9];	// matmul/matmul-hw.mlir:10996:16, :10997:12
  wire [31:0] _T_2688 = B_p0_rd_data[8'hEA];	// matmul/matmul-hw.mlir:10999:16, :11000:12
  wire [31:0] _T_2689 = B_p0_rd_data[8'hEB];	// matmul/matmul-hw.mlir:11002:16, :11003:12
  wire [31:0] _T_2690 = B_p0_rd_data[8'hEC];	// matmul/matmul-hw.mlir:11005:16, :11006:12
  wire [31:0] _T_2691 = B_p0_rd_data[8'hED];	// matmul/matmul-hw.mlir:11008:16, :11009:12
  wire [31:0] _T_2692 = B_p0_rd_data[8'hEE];	// matmul/matmul-hw.mlir:11011:16, :11012:12
  wire [31:0] _T_2693 = B_p0_rd_data[8'hEF];	// matmul/matmul-hw.mlir:11014:16, :11015:12
  wire [31:0] _T_2694 = B_p0_rd_data[8'hF0];	// matmul/matmul-hw.mlir:11017:16, :11018:12
  wire [31:0] _T_2695 = B_p0_rd_data[8'hF1];	// matmul/matmul-hw.mlir:11020:16, :11021:12
  wire [31:0] _T_2696 = B_p0_rd_data[8'hF2];	// matmul/matmul-hw.mlir:11023:16, :11024:12
  wire [31:0] _T_2697 = B_p0_rd_data[8'hF3];	// matmul/matmul-hw.mlir:11026:16, :11027:12
  wire [31:0] _T_2698 = B_p0_rd_data[8'hF4];	// matmul/matmul-hw.mlir:11029:16, :11030:12
  wire [31:0] _T_2699 = B_p0_rd_data[8'hF5];	// matmul/matmul-hw.mlir:11032:16, :11033:12
  wire [31:0] _T_2700 = B_p0_rd_data[8'hF6];	// matmul/matmul-hw.mlir:11035:16, :11036:12
  wire [31:0] _T_2701 = B_p0_rd_data[8'hF7];	// matmul/matmul-hw.mlir:11038:15, :11039:12
  wire [31:0] _T_2702 = B_p0_rd_data[8'hF8];	// matmul/matmul-hw.mlir:11041:15, :11042:12
  wire [31:0] _T_2703 = B_p0_rd_data[8'hF9];	// matmul/matmul-hw.mlir:11044:15, :11045:12
  wire [31:0] _T_2704 = B_p0_rd_data[8'hFA];	// matmul/matmul-hw.mlir:11047:15, :11048:12
  wire [31:0] _T_2705 = B_p0_rd_data[8'hFB];	// matmul/matmul-hw.mlir:11050:15, :11051:12
  wire [31:0] _T_2706 = B_p0_rd_data[8'hFC];	// matmul/matmul-hw.mlir:11053:15, :11054:12
  wire [31:0] _T_2707 = B_p0_rd_data[8'hFD];	// matmul/matmul-hw.mlir:11056:15, :11057:12
  wire [31:0] _T_2708 = B_p0_rd_data[8'hFE];	// matmul/matmul-hw.mlir:11059:15, :11060:12
  wire [31:0] _T_2709 = B_p0_rd_data[8'hFF];	// matmul/matmul-hw.mlir:11062:15, :11063:12
  localparam _T_2711 = 1'h0;	// matmul/matmul-hw.mlir:11146:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:11147:5
    if (rst)	// matmul/matmul-hw.mlir:11147:5
      _T_2710 <= _T_2711;	// matmul/matmul-hw.mlir:11150:7
    else	// matmul/matmul-hw.mlir:11147:5
      _T_2710 <= t;	// matmul/matmul-hw.mlir:11148:7
  end // always @(posedge)
  wire _T_2712 = _T_2710 & 1'h1 | _T_2189 & reg_1x1_r0_w1_inst3_p0_rd_data;	// matmul/matmul-hw.mlir:8029:13, :11145:12, :11155:12, :11156:12, :11157:12, :11178:39, :12484:12
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd6)
  ) reg_1x6_r0_w1_inst3 (	// matmul/matmul-hw.mlir:11167:39
    .p0_rd_en   (_T_2198),	// matmul/matmul-hw.mlir:11168:12
    .p1_wr_en   (_T_2197),	// matmul/matmul-hw.mlir:11171:12
    .p1_wr_data (_T_2196),	// matmul/matmul-hw.mlir:11172:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (reg_1x6_r0_w1_inst3_p0_rd_data)
  );
  assign _T_2198 = _T_2712 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :11168:12
  wire [5:0] _T_2713 = _T_2710 ? 6'h0 : reg_1x6_r0_w1_inst3_p0_rd_data;	// matmul/matmul-hw.mlir:8030:14, :11145:12, :11167:39, :11169:12
  wire [5:0] _T_2714 = _T_2713 + 6'h1;	// matmul/matmul-hw.mlir:8032:14, :11170:12
  assign _T_2197 = _T_2712 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :11171:12
  assign _T_2196 = _T_2712 ? _T_2714 : 6'bx;	// matmul/matmul-hw.mlir:10229:13, :11172:12
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd1)
  ) reg_1x1_r0_w1_inst3 (	// matmul/matmul-hw.mlir:11178:39
    .p0_rd_en   (_T_2193),	// matmul/matmul-hw.mlir:11181:12
    .p1_wr_en   (_T_2195),	// matmul/matmul-hw.mlir:11179:12
    .p1_wr_data (_T_2194),	// matmul/matmul-hw.mlir:11180:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (reg_1x1_r0_w1_inst3_p0_rd_data)
  );
  assign _T_2195 = _T_2712 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :11179:12
  assign _T_2194 = _T_2712 ? _T_2714 < 6'h10 : 1'bx;	// matmul/matmul-hw.mlir:8031:15, :10227:18, :11173:12, :11180:12
  assign _T_2193 = _T_2712 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :11181:12
  wire [4:0] _T_2715 = _T_2713[4:0];	// matmul/matmul-hw.mlir:11182:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:11184:5
    if (_T_2712)	// matmul/matmul-hw.mlir:11185:7
      _T_2716 <= _T_2715;	// matmul/matmul-hw.mlir:11186:9
  end // always @(posedge)
  wire [4:0] _T_2717 = _T_2712 ? _T_2715 : _T_2716;	// matmul/matmul-hw.mlir:11189:12, :11190:12
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank0 (	// matmul/matmul-hw.mlir:12215:31
    .p0_rd_en   (_T_2110),	// matmul/matmul-hw.mlir:13194:12
    .p1_wr_en   (_T_2187),	// matmul/matmul-hw.mlir:12491:12
    .p1_wr_data (_T_2186),	// matmul/matmul-hw.mlir:12492:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank0_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank1 (	// matmul/matmul-hw.mlir:12216:31
    .p0_rd_en   (_T_2107),	// matmul/matmul-hw.mlir:13197:12
    .p1_wr_en   (_T_2182),	// matmul/matmul-hw.mlir:12537:12
    .p1_wr_data (_T_2181),	// matmul/matmul-hw.mlir:12538:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank1_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank2 (	// matmul/matmul-hw.mlir:12217:31
    .p0_rd_en   (_T_2104),	// matmul/matmul-hw.mlir:13200:12
    .p1_wr_en   (_T_2177),	// matmul/matmul-hw.mlir:12583:12
    .p1_wr_data (_T_2176),	// matmul/matmul-hw.mlir:12584:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank2_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank3 (	// matmul/matmul-hw.mlir:12218:31
    .p0_rd_en   (_T_2101),	// matmul/matmul-hw.mlir:13203:12
    .p1_wr_en   (_T_2172),	// matmul/matmul-hw.mlir:12629:12
    .p1_wr_data (_T_2171),	// matmul/matmul-hw.mlir:12630:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank3_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank4 (	// matmul/matmul-hw.mlir:12219:31
    .p0_rd_en   (_T_2098),	// matmul/matmul-hw.mlir:13206:12
    .p1_wr_en   (_T_2167),	// matmul/matmul-hw.mlir:12675:12
    .p1_wr_data (_T_2166),	// matmul/matmul-hw.mlir:12676:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank4_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank5 (	// matmul/matmul-hw.mlir:12220:31
    .p0_rd_en   (_T_2095),	// matmul/matmul-hw.mlir:13209:12
    .p1_wr_en   (_T_2162),	// matmul/matmul-hw.mlir:12721:12
    .p1_wr_data (_T_2161),	// matmul/matmul-hw.mlir:12722:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank5_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank6 (	// matmul/matmul-hw.mlir:12221:31
    .p0_rd_en   (_T_2092),	// matmul/matmul-hw.mlir:13212:12
    .p1_wr_en   (_T_2157),	// matmul/matmul-hw.mlir:12767:12
    .p1_wr_data (_T_2156),	// matmul/matmul-hw.mlir:12768:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank6_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank7 (	// matmul/matmul-hw.mlir:12222:31
    .p0_rd_en   (_T_2089),	// matmul/matmul-hw.mlir:13215:12
    .p1_wr_en   (_T_2152),	// matmul/matmul-hw.mlir:12813:12
    .p1_wr_data (_T_2151),	// matmul/matmul-hw.mlir:12814:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank7_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank8 (	// matmul/matmul-hw.mlir:12223:31
    .p0_rd_en   (_T_2086),	// matmul/matmul-hw.mlir:13218:12
    .p1_wr_en   (_T_2147),	// matmul/matmul-hw.mlir:12859:12
    .p1_wr_data (_T_2146),	// matmul/matmul-hw.mlir:12860:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank8_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank9 (	// matmul/matmul-hw.mlir:12224:31
    .p0_rd_en   (_T_2083),	// matmul/matmul-hw.mlir:13221:12
    .p1_wr_en   (_T_2142),	// matmul/matmul-hw.mlir:12905:12
    .p1_wr_data (_T_2141),	// matmul/matmul-hw.mlir:12906:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank9_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank10 (	// matmul/matmul-hw.mlir:12225:32
    .p0_rd_en   (_T_2080),	// matmul/matmul-hw.mlir:13224:12
    .p1_wr_en   (_T_2137),	// matmul/matmul-hw.mlir:12951:12
    .p1_wr_data (_T_2136),	// matmul/matmul-hw.mlir:12952:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank10_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank11 (	// matmul/matmul-hw.mlir:12226:32
    .p0_rd_en   (_T_2077),	// matmul/matmul-hw.mlir:13227:12
    .p1_wr_en   (_T_2132),	// matmul/matmul-hw.mlir:12997:12
    .p1_wr_data (_T_2131),	// matmul/matmul-hw.mlir:12998:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank11_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank12 (	// matmul/matmul-hw.mlir:12227:32
    .p0_rd_en   (_T_2074),	// matmul/matmul-hw.mlir:13230:12
    .p1_wr_en   (_T_2127),	// matmul/matmul-hw.mlir:13043:12
    .p1_wr_data (_T_2126),	// matmul/matmul-hw.mlir:13044:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank12_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank13 (	// matmul/matmul-hw.mlir:12228:32
    .p0_rd_en   (_T_2071),	// matmul/matmul-hw.mlir:13233:12
    .p1_wr_en   (_T_2122),	// matmul/matmul-hw.mlir:13089:12
    .p1_wr_data (_T_2121),	// matmul/matmul-hw.mlir:13090:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank13_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank14 (	// matmul/matmul-hw.mlir:12229:32
    .p0_rd_en   (_T_2068),	// matmul/matmul-hw.mlir:13236:12
    .p1_wr_en   (_T_2117),	// matmul/matmul-hw.mlir:13135:12
    .p1_wr_data (_T_2116),	// matmul/matmul-hw.mlir:13136:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank14_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank15 (	// matmul/matmul-hw.mlir:12230:32
    .p0_rd_en   (_T_2065),	// matmul/matmul-hw.mlir:13254:12
    .p1_wr_en   (_T_2112),	// matmul/matmul-hw.mlir:13181:12
    .p1_wr_data (_T_2111),	// matmul/matmul-hw.mlir:13182:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank15_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank16 (	// matmul/matmul-hw.mlir:12231:32
    .p0_rd_en   (_T_2062),	// matmul/matmul-hw.mlir:13257:12
    .p1_wr_en   (_T_2109),	// matmul/matmul-hw.mlir:13195:12
    .p1_wr_data (_T_2108),	// matmul/matmul-hw.mlir:13196:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank16_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank17 (	// matmul/matmul-hw.mlir:12232:32
    .p0_rd_en   (_T_2059),	// matmul/matmul-hw.mlir:13260:12
    .p1_wr_en   (_T_2106),	// matmul/matmul-hw.mlir:13198:12
    .p1_wr_data (_T_2105),	// matmul/matmul-hw.mlir:13199:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank17_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank18 (	// matmul/matmul-hw.mlir:12233:32
    .p0_rd_en   (_T_2056),	// matmul/matmul-hw.mlir:13263:12
    .p1_wr_en   (_T_2103),	// matmul/matmul-hw.mlir:13201:12
    .p1_wr_data (_T_2102),	// matmul/matmul-hw.mlir:13202:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank18_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank19 (	// matmul/matmul-hw.mlir:12234:32
    .p0_rd_en   (_T_2053),	// matmul/matmul-hw.mlir:13266:12
    .p1_wr_en   (_T_2100),	// matmul/matmul-hw.mlir:13204:12
    .p1_wr_data (_T_2099),	// matmul/matmul-hw.mlir:13205:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank19_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank20 (	// matmul/matmul-hw.mlir:12235:32
    .p0_rd_en   (_T_2050),	// matmul/matmul-hw.mlir:13269:12
    .p1_wr_en   (_T_2097),	// matmul/matmul-hw.mlir:13207:12
    .p1_wr_data (_T_2096),	// matmul/matmul-hw.mlir:13208:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank20_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank21 (	// matmul/matmul-hw.mlir:12236:32
    .p0_rd_en   (_T_2047),	// matmul/matmul-hw.mlir:13272:12
    .p1_wr_en   (_T_2094),	// matmul/matmul-hw.mlir:13210:12
    .p1_wr_data (_T_2093),	// matmul/matmul-hw.mlir:13211:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank21_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank22 (	// matmul/matmul-hw.mlir:12237:32
    .p0_rd_en   (_T_2044),	// matmul/matmul-hw.mlir:13275:12
    .p1_wr_en   (_T_2091),	// matmul/matmul-hw.mlir:13213:12
    .p1_wr_data (_T_2090),	// matmul/matmul-hw.mlir:13214:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank22_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank23 (	// matmul/matmul-hw.mlir:12238:32
    .p0_rd_en   (_T_2041),	// matmul/matmul-hw.mlir:13278:12
    .p1_wr_en   (_T_2088),	// matmul/matmul-hw.mlir:13216:12
    .p1_wr_data (_T_2087),	// matmul/matmul-hw.mlir:13217:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank23_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank24 (	// matmul/matmul-hw.mlir:12239:32
    .p0_rd_en   (_T_2038),	// matmul/matmul-hw.mlir:13281:12
    .p1_wr_en   (_T_2085),	// matmul/matmul-hw.mlir:13219:12
    .p1_wr_data (_T_2084),	// matmul/matmul-hw.mlir:13220:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank24_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank25 (	// matmul/matmul-hw.mlir:12240:32
    .p0_rd_en   (_T_2035),	// matmul/matmul-hw.mlir:13284:12
    .p1_wr_en   (_T_2082),	// matmul/matmul-hw.mlir:13222:12
    .p1_wr_data (_T_2081),	// matmul/matmul-hw.mlir:13223:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank25_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank26 (	// matmul/matmul-hw.mlir:12241:32
    .p0_rd_en   (_T_2032),	// matmul/matmul-hw.mlir:13287:12
    .p1_wr_en   (_T_2079),	// matmul/matmul-hw.mlir:13225:12
    .p1_wr_data (_T_2078),	// matmul/matmul-hw.mlir:13226:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank26_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank27 (	// matmul/matmul-hw.mlir:12242:32
    .p0_rd_en   (_T_2029),	// matmul/matmul-hw.mlir:13290:12
    .p1_wr_en   (_T_2076),	// matmul/matmul-hw.mlir:13228:12
    .p1_wr_data (_T_2075),	// matmul/matmul-hw.mlir:13229:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank27_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank28 (	// matmul/matmul-hw.mlir:12243:32
    .p0_rd_en   (_T_2026),	// matmul/matmul-hw.mlir:13293:12
    .p1_wr_en   (_T_2073),	// matmul/matmul-hw.mlir:13231:12
    .p1_wr_data (_T_2072),	// matmul/matmul-hw.mlir:13232:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank28_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank29 (	// matmul/matmul-hw.mlir:12244:32
    .p0_rd_en   (_T_2023),	// matmul/matmul-hw.mlir:13296:12
    .p1_wr_en   (_T_2070),	// matmul/matmul-hw.mlir:13234:12
    .p1_wr_data (_T_2069),	// matmul/matmul-hw.mlir:13235:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank29_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank30 (	// matmul/matmul-hw.mlir:12245:32
    .p0_rd_en   (_T_2020),	// matmul/matmul-hw.mlir:13299:12
    .p1_wr_en   (_T_2067),	// matmul/matmul-hw.mlir:13237:12
    .p1_wr_data (_T_2066),	// matmul/matmul-hw.mlir:13238:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank30_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank31 (	// matmul/matmul-hw.mlir:12246:32
    .p0_rd_en   (_T_2017),	// matmul/matmul-hw.mlir:13317:12
    .p1_wr_en   (_T_2064),	// matmul/matmul-hw.mlir:13255:12
    .p1_wr_data (_T_2063),	// matmul/matmul-hw.mlir:13256:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank31_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank32 (	// matmul/matmul-hw.mlir:12247:32
    .p0_rd_en   (_T_2014),	// matmul/matmul-hw.mlir:13320:12
    .p1_wr_en   (_T_2061),	// matmul/matmul-hw.mlir:13258:12
    .p1_wr_data (_T_2060),	// matmul/matmul-hw.mlir:13259:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank32_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank33 (	// matmul/matmul-hw.mlir:12248:32
    .p0_rd_en   (_T_2011),	// matmul/matmul-hw.mlir:13323:12
    .p1_wr_en   (_T_2058),	// matmul/matmul-hw.mlir:13261:12
    .p1_wr_data (_T_2057),	// matmul/matmul-hw.mlir:13262:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank33_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank34 (	// matmul/matmul-hw.mlir:12249:32
    .p0_rd_en   (_T_2008),	// matmul/matmul-hw.mlir:13326:12
    .p1_wr_en   (_T_2055),	// matmul/matmul-hw.mlir:13264:12
    .p1_wr_data (_T_2054),	// matmul/matmul-hw.mlir:13265:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank34_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank35 (	// matmul/matmul-hw.mlir:12250:32
    .p0_rd_en   (_T_2005),	// matmul/matmul-hw.mlir:13329:12
    .p1_wr_en   (_T_2052),	// matmul/matmul-hw.mlir:13267:12
    .p1_wr_data (_T_2051),	// matmul/matmul-hw.mlir:13268:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank35_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank36 (	// matmul/matmul-hw.mlir:12251:32
    .p0_rd_en   (_T_2002),	// matmul/matmul-hw.mlir:13332:12
    .p1_wr_en   (_T_2049),	// matmul/matmul-hw.mlir:13270:12
    .p1_wr_data (_T_2048),	// matmul/matmul-hw.mlir:13271:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank36_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank37 (	// matmul/matmul-hw.mlir:12252:32
    .p0_rd_en   (_T_1999),	// matmul/matmul-hw.mlir:13335:12
    .p1_wr_en   (_T_2046),	// matmul/matmul-hw.mlir:13273:12
    .p1_wr_data (_T_2045),	// matmul/matmul-hw.mlir:13274:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank37_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank38 (	// matmul/matmul-hw.mlir:12253:32
    .p0_rd_en   (_T_1996),	// matmul/matmul-hw.mlir:13338:12
    .p1_wr_en   (_T_2043),	// matmul/matmul-hw.mlir:13276:12
    .p1_wr_data (_T_2042),	// matmul/matmul-hw.mlir:13277:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank38_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank39 (	// matmul/matmul-hw.mlir:12254:32
    .p0_rd_en   (_T_1993),	// matmul/matmul-hw.mlir:13341:12
    .p1_wr_en   (_T_2040),	// matmul/matmul-hw.mlir:13279:12
    .p1_wr_data (_T_2039),	// matmul/matmul-hw.mlir:13280:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank39_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank40 (	// matmul/matmul-hw.mlir:12255:32
    .p0_rd_en   (_T_1990),	// matmul/matmul-hw.mlir:13344:12
    .p1_wr_en   (_T_2037),	// matmul/matmul-hw.mlir:13282:12
    .p1_wr_data (_T_2036),	// matmul/matmul-hw.mlir:13283:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank40_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank41 (	// matmul/matmul-hw.mlir:12256:32
    .p0_rd_en   (_T_1987),	// matmul/matmul-hw.mlir:13347:12
    .p1_wr_en   (_T_2034),	// matmul/matmul-hw.mlir:13285:12
    .p1_wr_data (_T_2033),	// matmul/matmul-hw.mlir:13286:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank41_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank42 (	// matmul/matmul-hw.mlir:12257:32
    .p0_rd_en   (_T_1984),	// matmul/matmul-hw.mlir:13350:12
    .p1_wr_en   (_T_2031),	// matmul/matmul-hw.mlir:13288:12
    .p1_wr_data (_T_2030),	// matmul/matmul-hw.mlir:13289:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank42_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank43 (	// matmul/matmul-hw.mlir:12258:32
    .p0_rd_en   (_T_1981),	// matmul/matmul-hw.mlir:13353:12
    .p1_wr_en   (_T_2028),	// matmul/matmul-hw.mlir:13291:12
    .p1_wr_data (_T_2027),	// matmul/matmul-hw.mlir:13292:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank43_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank44 (	// matmul/matmul-hw.mlir:12259:32
    .p0_rd_en   (_T_1978),	// matmul/matmul-hw.mlir:13356:12
    .p1_wr_en   (_T_2025),	// matmul/matmul-hw.mlir:13294:12
    .p1_wr_data (_T_2024),	// matmul/matmul-hw.mlir:13295:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank44_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank45 (	// matmul/matmul-hw.mlir:12260:32
    .p0_rd_en   (_T_1975),	// matmul/matmul-hw.mlir:13359:12
    .p1_wr_en   (_T_2022),	// matmul/matmul-hw.mlir:13297:12
    .p1_wr_data (_T_2021),	// matmul/matmul-hw.mlir:13298:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank45_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank46 (	// matmul/matmul-hw.mlir:12261:32
    .p0_rd_en   (_T_1972),	// matmul/matmul-hw.mlir:13362:12
    .p1_wr_en   (_T_2019),	// matmul/matmul-hw.mlir:13300:12
    .p1_wr_data (_T_2018),	// matmul/matmul-hw.mlir:13301:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank46_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank47 (	// matmul/matmul-hw.mlir:12262:32
    .p0_rd_en   (_T_1969),	// matmul/matmul-hw.mlir:13380:12
    .p1_wr_en   (_T_2016),	// matmul/matmul-hw.mlir:13318:12
    .p1_wr_data (_T_2015),	// matmul/matmul-hw.mlir:13319:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank47_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank48 (	// matmul/matmul-hw.mlir:12263:32
    .p0_rd_en   (_T_1966),	// matmul/matmul-hw.mlir:13383:12
    .p1_wr_en   (_T_2013),	// matmul/matmul-hw.mlir:13321:12
    .p1_wr_data (_T_2012),	// matmul/matmul-hw.mlir:13322:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank48_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank49 (	// matmul/matmul-hw.mlir:12264:32
    .p0_rd_en   (_T_1963),	// matmul/matmul-hw.mlir:13386:12
    .p1_wr_en   (_T_2010),	// matmul/matmul-hw.mlir:13324:12
    .p1_wr_data (_T_2009),	// matmul/matmul-hw.mlir:13325:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank49_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank50 (	// matmul/matmul-hw.mlir:12265:32
    .p0_rd_en   (_T_1960),	// matmul/matmul-hw.mlir:13389:12
    .p1_wr_en   (_T_2007),	// matmul/matmul-hw.mlir:13327:12
    .p1_wr_data (_T_2006),	// matmul/matmul-hw.mlir:13328:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank50_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank51 (	// matmul/matmul-hw.mlir:12266:32
    .p0_rd_en   (_T_1957),	// matmul/matmul-hw.mlir:13392:12
    .p1_wr_en   (_T_2004),	// matmul/matmul-hw.mlir:13330:12
    .p1_wr_data (_T_2003),	// matmul/matmul-hw.mlir:13331:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank51_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank52 (	// matmul/matmul-hw.mlir:12267:32
    .p0_rd_en   (_T_1954),	// matmul/matmul-hw.mlir:13395:12
    .p1_wr_en   (_T_2001),	// matmul/matmul-hw.mlir:13333:12
    .p1_wr_data (_T_2000),	// matmul/matmul-hw.mlir:13334:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank52_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank53 (	// matmul/matmul-hw.mlir:12268:32
    .p0_rd_en   (_T_1951),	// matmul/matmul-hw.mlir:13398:12
    .p1_wr_en   (_T_1998),	// matmul/matmul-hw.mlir:13336:12
    .p1_wr_data (_T_1997),	// matmul/matmul-hw.mlir:13337:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank53_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank54 (	// matmul/matmul-hw.mlir:12269:32
    .p0_rd_en   (_T_1948),	// matmul/matmul-hw.mlir:13401:12
    .p1_wr_en   (_T_1995),	// matmul/matmul-hw.mlir:13339:12
    .p1_wr_data (_T_1994),	// matmul/matmul-hw.mlir:13340:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank54_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank55 (	// matmul/matmul-hw.mlir:12270:32
    .p0_rd_en   (_T_1945),	// matmul/matmul-hw.mlir:13404:12
    .p1_wr_en   (_T_1992),	// matmul/matmul-hw.mlir:13342:12
    .p1_wr_data (_T_1991),	// matmul/matmul-hw.mlir:13343:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank55_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank56 (	// matmul/matmul-hw.mlir:12271:32
    .p0_rd_en   (_T_1942),	// matmul/matmul-hw.mlir:13407:12
    .p1_wr_en   (_T_1989),	// matmul/matmul-hw.mlir:13345:12
    .p1_wr_data (_T_1988),	// matmul/matmul-hw.mlir:13346:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank56_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank57 (	// matmul/matmul-hw.mlir:12272:32
    .p0_rd_en   (_T_1939),	// matmul/matmul-hw.mlir:13410:12
    .p1_wr_en   (_T_1986),	// matmul/matmul-hw.mlir:13348:12
    .p1_wr_data (_T_1985),	// matmul/matmul-hw.mlir:13349:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank57_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank58 (	// matmul/matmul-hw.mlir:12273:32
    .p0_rd_en   (_T_1936),	// matmul/matmul-hw.mlir:13413:12
    .p1_wr_en   (_T_1983),	// matmul/matmul-hw.mlir:13351:12
    .p1_wr_data (_T_1982),	// matmul/matmul-hw.mlir:13352:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank58_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank59 (	// matmul/matmul-hw.mlir:12274:32
    .p0_rd_en   (_T_1933),	// matmul/matmul-hw.mlir:13416:12
    .p1_wr_en   (_T_1980),	// matmul/matmul-hw.mlir:13354:12
    .p1_wr_data (_T_1979),	// matmul/matmul-hw.mlir:13355:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank59_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank60 (	// matmul/matmul-hw.mlir:12275:32
    .p0_rd_en   (_T_1930),	// matmul/matmul-hw.mlir:13419:12
    .p1_wr_en   (_T_1977),	// matmul/matmul-hw.mlir:13357:12
    .p1_wr_data (_T_1976),	// matmul/matmul-hw.mlir:13358:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank60_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank61 (	// matmul/matmul-hw.mlir:12276:32
    .p0_rd_en   (_T_1927),	// matmul/matmul-hw.mlir:13422:12
    .p1_wr_en   (_T_1974),	// matmul/matmul-hw.mlir:13360:12
    .p1_wr_data (_T_1973),	// matmul/matmul-hw.mlir:13361:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank61_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank62 (	// matmul/matmul-hw.mlir:12277:32
    .p0_rd_en   (_T_1924),	// matmul/matmul-hw.mlir:13425:12
    .p1_wr_en   (_T_1971),	// matmul/matmul-hw.mlir:13363:12
    .p1_wr_data (_T_1970),	// matmul/matmul-hw.mlir:13364:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank62_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank63 (	// matmul/matmul-hw.mlir:12278:32
    .p0_rd_en   (_T_1921),	// matmul/matmul-hw.mlir:13443:12
    .p1_wr_en   (_T_1968),	// matmul/matmul-hw.mlir:13381:12
    .p1_wr_data (_T_1967),	// matmul/matmul-hw.mlir:13382:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank63_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank64 (	// matmul/matmul-hw.mlir:12279:32
    .p0_rd_en   (_T_1918),	// matmul/matmul-hw.mlir:13446:12
    .p1_wr_en   (_T_1965),	// matmul/matmul-hw.mlir:13384:12
    .p1_wr_data (_T_1964),	// matmul/matmul-hw.mlir:13385:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank64_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank65 (	// matmul/matmul-hw.mlir:12280:32
    .p0_rd_en   (_T_1915),	// matmul/matmul-hw.mlir:13449:12
    .p1_wr_en   (_T_1962),	// matmul/matmul-hw.mlir:13387:12
    .p1_wr_data (_T_1961),	// matmul/matmul-hw.mlir:13388:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank65_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank66 (	// matmul/matmul-hw.mlir:12281:32
    .p0_rd_en   (_T_1912),	// matmul/matmul-hw.mlir:13452:12
    .p1_wr_en   (_T_1959),	// matmul/matmul-hw.mlir:13390:12
    .p1_wr_data (_T_1958),	// matmul/matmul-hw.mlir:13391:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank66_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank67 (	// matmul/matmul-hw.mlir:12282:32
    .p0_rd_en   (_T_1909),	// matmul/matmul-hw.mlir:13455:12
    .p1_wr_en   (_T_1956),	// matmul/matmul-hw.mlir:13393:12
    .p1_wr_data (_T_1955),	// matmul/matmul-hw.mlir:13394:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank67_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank68 (	// matmul/matmul-hw.mlir:12283:32
    .p0_rd_en   (_T_1906),	// matmul/matmul-hw.mlir:13458:12
    .p1_wr_en   (_T_1953),	// matmul/matmul-hw.mlir:13396:12
    .p1_wr_data (_T_1952),	// matmul/matmul-hw.mlir:13397:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank68_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank69 (	// matmul/matmul-hw.mlir:12284:32
    .p0_rd_en   (_T_1903),	// matmul/matmul-hw.mlir:13461:12
    .p1_wr_en   (_T_1950),	// matmul/matmul-hw.mlir:13399:12
    .p1_wr_data (_T_1949),	// matmul/matmul-hw.mlir:13400:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank69_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank70 (	// matmul/matmul-hw.mlir:12285:32
    .p0_rd_en   (_T_1900),	// matmul/matmul-hw.mlir:13464:12
    .p1_wr_en   (_T_1947),	// matmul/matmul-hw.mlir:13402:12
    .p1_wr_data (_T_1946),	// matmul/matmul-hw.mlir:13403:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank70_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank71 (	// matmul/matmul-hw.mlir:12286:32
    .p0_rd_en   (_T_1897),	// matmul/matmul-hw.mlir:13467:12
    .p1_wr_en   (_T_1944),	// matmul/matmul-hw.mlir:13405:12
    .p1_wr_data (_T_1943),	// matmul/matmul-hw.mlir:13406:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank71_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank72 (	// matmul/matmul-hw.mlir:12287:32
    .p0_rd_en   (_T_1894),	// matmul/matmul-hw.mlir:13470:12
    .p1_wr_en   (_T_1941),	// matmul/matmul-hw.mlir:13408:12
    .p1_wr_data (_T_1940),	// matmul/matmul-hw.mlir:13409:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank72_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank73 (	// matmul/matmul-hw.mlir:12288:32
    .p0_rd_en   (_T_1891),	// matmul/matmul-hw.mlir:13473:12
    .p1_wr_en   (_T_1938),	// matmul/matmul-hw.mlir:13411:12
    .p1_wr_data (_T_1937),	// matmul/matmul-hw.mlir:13412:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank73_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank74 (	// matmul/matmul-hw.mlir:12289:32
    .p0_rd_en   (_T_1888),	// matmul/matmul-hw.mlir:13476:12
    .p1_wr_en   (_T_1935),	// matmul/matmul-hw.mlir:13414:12
    .p1_wr_data (_T_1934),	// matmul/matmul-hw.mlir:13415:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank74_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank75 (	// matmul/matmul-hw.mlir:12290:32
    .p0_rd_en   (_T_1885),	// matmul/matmul-hw.mlir:13479:12
    .p1_wr_en   (_T_1932),	// matmul/matmul-hw.mlir:13417:12
    .p1_wr_data (_T_1931),	// matmul/matmul-hw.mlir:13418:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank75_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank76 (	// matmul/matmul-hw.mlir:12291:32
    .p0_rd_en   (_T_1882),	// matmul/matmul-hw.mlir:13482:12
    .p1_wr_en   (_T_1929),	// matmul/matmul-hw.mlir:13420:12
    .p1_wr_data (_T_1928),	// matmul/matmul-hw.mlir:13421:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank76_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank77 (	// matmul/matmul-hw.mlir:12292:32
    .p0_rd_en   (_T_1879),	// matmul/matmul-hw.mlir:13485:12
    .p1_wr_en   (_T_1926),	// matmul/matmul-hw.mlir:13423:12
    .p1_wr_data (_T_1925),	// matmul/matmul-hw.mlir:13424:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank77_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank78 (	// matmul/matmul-hw.mlir:12293:32
    .p0_rd_en   (_T_1876),	// matmul/matmul-hw.mlir:13488:12
    .p1_wr_en   (_T_1923),	// matmul/matmul-hw.mlir:13426:12
    .p1_wr_data (_T_1922),	// matmul/matmul-hw.mlir:13427:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank78_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank79 (	// matmul/matmul-hw.mlir:12294:32
    .p0_rd_en   (_T_1873),	// matmul/matmul-hw.mlir:13506:12
    .p1_wr_en   (_T_1920),	// matmul/matmul-hw.mlir:13444:12
    .p1_wr_data (_T_1919),	// matmul/matmul-hw.mlir:13445:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank79_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank80 (	// matmul/matmul-hw.mlir:12295:32
    .p0_rd_en   (_T_1870),	// matmul/matmul-hw.mlir:13509:12
    .p1_wr_en   (_T_1917),	// matmul/matmul-hw.mlir:13447:12
    .p1_wr_data (_T_1916),	// matmul/matmul-hw.mlir:13448:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank80_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank81 (	// matmul/matmul-hw.mlir:12296:32
    .p0_rd_en   (_T_1867),	// matmul/matmul-hw.mlir:13512:12
    .p1_wr_en   (_T_1914),	// matmul/matmul-hw.mlir:13450:12
    .p1_wr_data (_T_1913),	// matmul/matmul-hw.mlir:13451:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank81_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank82 (	// matmul/matmul-hw.mlir:12297:32
    .p0_rd_en   (_T_1864),	// matmul/matmul-hw.mlir:13515:12
    .p1_wr_en   (_T_1911),	// matmul/matmul-hw.mlir:13453:12
    .p1_wr_data (_T_1910),	// matmul/matmul-hw.mlir:13454:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank82_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank83 (	// matmul/matmul-hw.mlir:12298:32
    .p0_rd_en   (_T_1861),	// matmul/matmul-hw.mlir:13518:12
    .p1_wr_en   (_T_1908),	// matmul/matmul-hw.mlir:13456:12
    .p1_wr_data (_T_1907),	// matmul/matmul-hw.mlir:13457:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank83_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank84 (	// matmul/matmul-hw.mlir:12299:32
    .p0_rd_en   (_T_1858),	// matmul/matmul-hw.mlir:13521:12
    .p1_wr_en   (_T_1905),	// matmul/matmul-hw.mlir:13459:12
    .p1_wr_data (_T_1904),	// matmul/matmul-hw.mlir:13460:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank84_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank85 (	// matmul/matmul-hw.mlir:12300:32
    .p0_rd_en   (_T_1855),	// matmul/matmul-hw.mlir:13524:12
    .p1_wr_en   (_T_1902),	// matmul/matmul-hw.mlir:13462:12
    .p1_wr_data (_T_1901),	// matmul/matmul-hw.mlir:13463:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank85_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank86 (	// matmul/matmul-hw.mlir:12301:32
    .p0_rd_en   (_T_1852),	// matmul/matmul-hw.mlir:13527:12
    .p1_wr_en   (_T_1899),	// matmul/matmul-hw.mlir:13465:12
    .p1_wr_data (_T_1898),	// matmul/matmul-hw.mlir:13466:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank86_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank87 (	// matmul/matmul-hw.mlir:12302:32
    .p0_rd_en   (_T_1849),	// matmul/matmul-hw.mlir:13530:12
    .p1_wr_en   (_T_1896),	// matmul/matmul-hw.mlir:13468:12
    .p1_wr_data (_T_1895),	// matmul/matmul-hw.mlir:13469:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank87_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank88 (	// matmul/matmul-hw.mlir:12303:32
    .p0_rd_en   (_T_1846),	// matmul/matmul-hw.mlir:13533:12
    .p1_wr_en   (_T_1893),	// matmul/matmul-hw.mlir:13471:12
    .p1_wr_data (_T_1892),	// matmul/matmul-hw.mlir:13472:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank88_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank89 (	// matmul/matmul-hw.mlir:12304:32
    .p0_rd_en   (_T_1843),	// matmul/matmul-hw.mlir:13536:12
    .p1_wr_en   (_T_1890),	// matmul/matmul-hw.mlir:13474:12
    .p1_wr_data (_T_1889),	// matmul/matmul-hw.mlir:13475:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank89_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank90 (	// matmul/matmul-hw.mlir:12305:32
    .p0_rd_en   (_T_1840),	// matmul/matmul-hw.mlir:13539:12
    .p1_wr_en   (_T_1887),	// matmul/matmul-hw.mlir:13477:12
    .p1_wr_data (_T_1886),	// matmul/matmul-hw.mlir:13478:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank90_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank91 (	// matmul/matmul-hw.mlir:12306:32
    .p0_rd_en   (_T_1837),	// matmul/matmul-hw.mlir:13542:12
    .p1_wr_en   (_T_1884),	// matmul/matmul-hw.mlir:13480:12
    .p1_wr_data (_T_1883),	// matmul/matmul-hw.mlir:13481:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank91_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank92 (	// matmul/matmul-hw.mlir:12307:32
    .p0_rd_en   (_T_1834),	// matmul/matmul-hw.mlir:13545:12
    .p1_wr_en   (_T_1881),	// matmul/matmul-hw.mlir:13483:12
    .p1_wr_data (_T_1880),	// matmul/matmul-hw.mlir:13484:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank92_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank93 (	// matmul/matmul-hw.mlir:12308:32
    .p0_rd_en   (_T_1831),	// matmul/matmul-hw.mlir:13548:12
    .p1_wr_en   (_T_1878),	// matmul/matmul-hw.mlir:13486:12
    .p1_wr_data (_T_1877),	// matmul/matmul-hw.mlir:13487:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank93_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank94 (	// matmul/matmul-hw.mlir:12309:32
    .p0_rd_en   (_T_1828),	// matmul/matmul-hw.mlir:13551:12
    .p1_wr_en   (_T_1875),	// matmul/matmul-hw.mlir:13489:12
    .p1_wr_data (_T_1874),	// matmul/matmul-hw.mlir:13490:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank94_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank95 (	// matmul/matmul-hw.mlir:12310:32
    .p0_rd_en   (_T_1825),	// matmul/matmul-hw.mlir:13569:12
    .p1_wr_en   (_T_1872),	// matmul/matmul-hw.mlir:13507:12
    .p1_wr_data (_T_1871),	// matmul/matmul-hw.mlir:13508:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank95_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank96 (	// matmul/matmul-hw.mlir:12311:32
    .p0_rd_en   (_T_1822),	// matmul/matmul-hw.mlir:13572:12
    .p1_wr_en   (_T_1869),	// matmul/matmul-hw.mlir:13510:12
    .p1_wr_data (_T_1868),	// matmul/matmul-hw.mlir:13511:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank96_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank97 (	// matmul/matmul-hw.mlir:12312:32
    .p0_rd_en   (_T_1819),	// matmul/matmul-hw.mlir:13575:12
    .p1_wr_en   (_T_1866),	// matmul/matmul-hw.mlir:13513:12
    .p1_wr_data (_T_1865),	// matmul/matmul-hw.mlir:13514:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank97_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank98 (	// matmul/matmul-hw.mlir:12313:32
    .p0_rd_en   (_T_1816),	// matmul/matmul-hw.mlir:13578:12
    .p1_wr_en   (_T_1863),	// matmul/matmul-hw.mlir:13516:12
    .p1_wr_data (_T_1862),	// matmul/matmul-hw.mlir:13517:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank98_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank99 (	// matmul/matmul-hw.mlir:12314:32
    .p0_rd_en   (_T_1813),	// matmul/matmul-hw.mlir:13581:12
    .p1_wr_en   (_T_1860),	// matmul/matmul-hw.mlir:13519:12
    .p1_wr_data (_T_1859),	// matmul/matmul-hw.mlir:13520:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank99_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank100 (	// matmul/matmul-hw.mlir:12315:33
    .p0_rd_en   (_T_1810),	// matmul/matmul-hw.mlir:13584:12
    .p1_wr_en   (_T_1857),	// matmul/matmul-hw.mlir:13522:12
    .p1_wr_data (_T_1856),	// matmul/matmul-hw.mlir:13523:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank100_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank101 (	// matmul/matmul-hw.mlir:12316:33
    .p0_rd_en   (_T_1807),	// matmul/matmul-hw.mlir:13587:12
    .p1_wr_en   (_T_1854),	// matmul/matmul-hw.mlir:13525:12
    .p1_wr_data (_T_1853),	// matmul/matmul-hw.mlir:13526:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank101_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank102 (	// matmul/matmul-hw.mlir:12317:33
    .p0_rd_en   (_T_1804),	// matmul/matmul-hw.mlir:13590:12
    .p1_wr_en   (_T_1851),	// matmul/matmul-hw.mlir:13528:12
    .p1_wr_data (_T_1850),	// matmul/matmul-hw.mlir:13529:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank102_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank103 (	// matmul/matmul-hw.mlir:12318:33
    .p0_rd_en   (_T_1801),	// matmul/matmul-hw.mlir:13593:12
    .p1_wr_en   (_T_1848),	// matmul/matmul-hw.mlir:13531:12
    .p1_wr_data (_T_1847),	// matmul/matmul-hw.mlir:13532:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank103_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank104 (	// matmul/matmul-hw.mlir:12319:33
    .p0_rd_en   (_T_1798),	// matmul/matmul-hw.mlir:13596:12
    .p1_wr_en   (_T_1845),	// matmul/matmul-hw.mlir:13534:12
    .p1_wr_data (_T_1844),	// matmul/matmul-hw.mlir:13535:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank104_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank105 (	// matmul/matmul-hw.mlir:12320:33
    .p0_rd_en   (_T_1795),	// matmul/matmul-hw.mlir:13599:12
    .p1_wr_en   (_T_1842),	// matmul/matmul-hw.mlir:13537:12
    .p1_wr_data (_T_1841),	// matmul/matmul-hw.mlir:13538:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank105_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank106 (	// matmul/matmul-hw.mlir:12321:33
    .p0_rd_en   (_T_1792),	// matmul/matmul-hw.mlir:13602:12
    .p1_wr_en   (_T_1839),	// matmul/matmul-hw.mlir:13540:12
    .p1_wr_data (_T_1838),	// matmul/matmul-hw.mlir:13541:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank106_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank107 (	// matmul/matmul-hw.mlir:12322:33
    .p0_rd_en   (_T_1789),	// matmul/matmul-hw.mlir:13605:12
    .p1_wr_en   (_T_1836),	// matmul/matmul-hw.mlir:13543:12
    .p1_wr_data (_T_1835),	// matmul/matmul-hw.mlir:13544:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank107_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank108 (	// matmul/matmul-hw.mlir:12323:33
    .p0_rd_en   (_T_1786),	// matmul/matmul-hw.mlir:13608:12
    .p1_wr_en   (_T_1833),	// matmul/matmul-hw.mlir:13546:12
    .p1_wr_data (_T_1832),	// matmul/matmul-hw.mlir:13547:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank108_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank109 (	// matmul/matmul-hw.mlir:12324:33
    .p0_rd_en   (_T_1783),	// matmul/matmul-hw.mlir:13611:12
    .p1_wr_en   (_T_1830),	// matmul/matmul-hw.mlir:13549:12
    .p1_wr_data (_T_1829),	// matmul/matmul-hw.mlir:13550:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank109_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank110 (	// matmul/matmul-hw.mlir:12325:33
    .p0_rd_en   (_T_1780),	// matmul/matmul-hw.mlir:13614:12
    .p1_wr_en   (_T_1827),	// matmul/matmul-hw.mlir:13552:12
    .p1_wr_data (_T_1826),	// matmul/matmul-hw.mlir:13553:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank110_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank111 (	// matmul/matmul-hw.mlir:12326:33
    .p0_rd_en   (_T_1777),	// matmul/matmul-hw.mlir:13632:12
    .p1_wr_en   (_T_1824),	// matmul/matmul-hw.mlir:13570:12
    .p1_wr_data (_T_1823),	// matmul/matmul-hw.mlir:13571:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank111_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank112 (	// matmul/matmul-hw.mlir:12327:33
    .p0_rd_en   (_T_1774),	// matmul/matmul-hw.mlir:13635:12
    .p1_wr_en   (_T_1821),	// matmul/matmul-hw.mlir:13573:12
    .p1_wr_data (_T_1820),	// matmul/matmul-hw.mlir:13574:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank112_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank113 (	// matmul/matmul-hw.mlir:12328:33
    .p0_rd_en   (_T_1771),	// matmul/matmul-hw.mlir:13638:13
    .p1_wr_en   (_T_1818),	// matmul/matmul-hw.mlir:13576:12
    .p1_wr_data (_T_1817),	// matmul/matmul-hw.mlir:13577:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank113_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank114 (	// matmul/matmul-hw.mlir:12329:33
    .p0_rd_en   (_T_1768),	// matmul/matmul-hw.mlir:13641:13
    .p1_wr_en   (_T_1815),	// matmul/matmul-hw.mlir:13579:12
    .p1_wr_data (_T_1814),	// matmul/matmul-hw.mlir:13580:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank114_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank115 (	// matmul/matmul-hw.mlir:12330:33
    .p0_rd_en   (_T_1765),	// matmul/matmul-hw.mlir:13644:13
    .p1_wr_en   (_T_1812),	// matmul/matmul-hw.mlir:13582:12
    .p1_wr_data (_T_1811),	// matmul/matmul-hw.mlir:13583:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank115_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank116 (	// matmul/matmul-hw.mlir:12331:33
    .p0_rd_en   (_T_1762),	// matmul/matmul-hw.mlir:13647:13
    .p1_wr_en   (_T_1809),	// matmul/matmul-hw.mlir:13585:12
    .p1_wr_data (_T_1808),	// matmul/matmul-hw.mlir:13586:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank116_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank117 (	// matmul/matmul-hw.mlir:12332:33
    .p0_rd_en   (_T_1759),	// matmul/matmul-hw.mlir:13650:13
    .p1_wr_en   (_T_1806),	// matmul/matmul-hw.mlir:13588:12
    .p1_wr_data (_T_1805),	// matmul/matmul-hw.mlir:13589:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank117_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank118 (	// matmul/matmul-hw.mlir:12333:33
    .p0_rd_en   (_T_1756),	// matmul/matmul-hw.mlir:13653:13
    .p1_wr_en   (_T_1803),	// matmul/matmul-hw.mlir:13591:12
    .p1_wr_data (_T_1802),	// matmul/matmul-hw.mlir:13592:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank118_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank119 (	// matmul/matmul-hw.mlir:12334:33
    .p0_rd_en   (_T_1753),	// matmul/matmul-hw.mlir:13656:13
    .p1_wr_en   (_T_1800),	// matmul/matmul-hw.mlir:13594:12
    .p1_wr_data (_T_1799),	// matmul/matmul-hw.mlir:13595:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank119_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank120 (	// matmul/matmul-hw.mlir:12335:33
    .p0_rd_en   (_T_1750),	// matmul/matmul-hw.mlir:13659:13
    .p1_wr_en   (_T_1797),	// matmul/matmul-hw.mlir:13597:12
    .p1_wr_data (_T_1796),	// matmul/matmul-hw.mlir:13598:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank120_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank121 (	// matmul/matmul-hw.mlir:12336:33
    .p0_rd_en   (_T_1747),	// matmul/matmul-hw.mlir:13662:13
    .p1_wr_en   (_T_1794),	// matmul/matmul-hw.mlir:13600:12
    .p1_wr_data (_T_1793),	// matmul/matmul-hw.mlir:13601:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank121_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank122 (	// matmul/matmul-hw.mlir:12337:33
    .p0_rd_en   (_T_1744),	// matmul/matmul-hw.mlir:13665:13
    .p1_wr_en   (_T_1791),	// matmul/matmul-hw.mlir:13603:12
    .p1_wr_data (_T_1790),	// matmul/matmul-hw.mlir:13604:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank122_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank123 (	// matmul/matmul-hw.mlir:12338:33
    .p0_rd_en   (_T_1741),	// matmul/matmul-hw.mlir:13668:13
    .p1_wr_en   (_T_1788),	// matmul/matmul-hw.mlir:13606:12
    .p1_wr_data (_T_1787),	// matmul/matmul-hw.mlir:13607:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank123_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank124 (	// matmul/matmul-hw.mlir:12339:33
    .p0_rd_en   (_T_1738),	// matmul/matmul-hw.mlir:13671:13
    .p1_wr_en   (_T_1785),	// matmul/matmul-hw.mlir:13609:12
    .p1_wr_data (_T_1784),	// matmul/matmul-hw.mlir:13610:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank124_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank125 (	// matmul/matmul-hw.mlir:12340:33
    .p0_rd_en   (_T_1735),	// matmul/matmul-hw.mlir:13674:13
    .p1_wr_en   (_T_1782),	// matmul/matmul-hw.mlir:13612:12
    .p1_wr_data (_T_1781),	// matmul/matmul-hw.mlir:13613:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank125_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank126 (	// matmul/matmul-hw.mlir:12341:33
    .p0_rd_en   (_T_1732),	// matmul/matmul-hw.mlir:13677:13
    .p1_wr_en   (_T_1779),	// matmul/matmul-hw.mlir:13615:12
    .p1_wr_data (_T_1778),	// matmul/matmul-hw.mlir:13616:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank126_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank127 (	// matmul/matmul-hw.mlir:12342:33
    .p0_rd_en   (_T_1729),	// matmul/matmul-hw.mlir:13695:13
    .p1_wr_en   (_T_1776),	// matmul/matmul-hw.mlir:13633:12
    .p1_wr_data (_T_1775),	// matmul/matmul-hw.mlir:13634:12
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank127_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank128 (	// matmul/matmul-hw.mlir:12343:33
    .p0_rd_en   (_T_1726),	// matmul/matmul-hw.mlir:13698:13
    .p1_wr_en   (_T_1773),	// matmul/matmul-hw.mlir:13636:13
    .p1_wr_data (_T_1772),	// matmul/matmul-hw.mlir:13637:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank128_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank129 (	// matmul/matmul-hw.mlir:12344:33
    .p0_rd_en   (_T_1723),	// matmul/matmul-hw.mlir:13701:13
    .p1_wr_en   (_T_1770),	// matmul/matmul-hw.mlir:13639:13
    .p1_wr_data (_T_1769),	// matmul/matmul-hw.mlir:13640:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank129_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank130 (	// matmul/matmul-hw.mlir:12345:33
    .p0_rd_en   (_T_1720),	// matmul/matmul-hw.mlir:13704:13
    .p1_wr_en   (_T_1767),	// matmul/matmul-hw.mlir:13642:13
    .p1_wr_data (_T_1766),	// matmul/matmul-hw.mlir:13643:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank130_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank131 (	// matmul/matmul-hw.mlir:12346:33
    .p0_rd_en   (_T_1717),	// matmul/matmul-hw.mlir:13707:13
    .p1_wr_en   (_T_1764),	// matmul/matmul-hw.mlir:13645:13
    .p1_wr_data (_T_1763),	// matmul/matmul-hw.mlir:13646:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank131_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank132 (	// matmul/matmul-hw.mlir:12347:33
    .p0_rd_en   (_T_1714),	// matmul/matmul-hw.mlir:13710:13
    .p1_wr_en   (_T_1761),	// matmul/matmul-hw.mlir:13648:13
    .p1_wr_data (_T_1760),	// matmul/matmul-hw.mlir:13649:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank132_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank133 (	// matmul/matmul-hw.mlir:12348:33
    .p0_rd_en   (_T_1711),	// matmul/matmul-hw.mlir:13713:13
    .p1_wr_en   (_T_1758),	// matmul/matmul-hw.mlir:13651:13
    .p1_wr_data (_T_1757),	// matmul/matmul-hw.mlir:13652:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank133_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank134 (	// matmul/matmul-hw.mlir:12349:33
    .p0_rd_en   (_T_1708),	// matmul/matmul-hw.mlir:13716:13
    .p1_wr_en   (_T_1755),	// matmul/matmul-hw.mlir:13654:13
    .p1_wr_data (_T_1754),	// matmul/matmul-hw.mlir:13655:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank134_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank135 (	// matmul/matmul-hw.mlir:12350:33
    .p0_rd_en   (_T_1705),	// matmul/matmul-hw.mlir:13719:13
    .p1_wr_en   (_T_1752),	// matmul/matmul-hw.mlir:13657:13
    .p1_wr_data (_T_1751),	// matmul/matmul-hw.mlir:13658:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank135_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank136 (	// matmul/matmul-hw.mlir:12351:33
    .p0_rd_en   (_T_1702),	// matmul/matmul-hw.mlir:13722:13
    .p1_wr_en   (_T_1749),	// matmul/matmul-hw.mlir:13660:13
    .p1_wr_data (_T_1748),	// matmul/matmul-hw.mlir:13661:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank136_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank137 (	// matmul/matmul-hw.mlir:12352:33
    .p0_rd_en   (_T_1699),	// matmul/matmul-hw.mlir:13725:13
    .p1_wr_en   (_T_1746),	// matmul/matmul-hw.mlir:13663:13
    .p1_wr_data (_T_1745),	// matmul/matmul-hw.mlir:13664:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank137_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank138 (	// matmul/matmul-hw.mlir:12353:33
    .p0_rd_en   (_T_1696),	// matmul/matmul-hw.mlir:13728:13
    .p1_wr_en   (_T_1743),	// matmul/matmul-hw.mlir:13666:13
    .p1_wr_data (_T_1742),	// matmul/matmul-hw.mlir:13667:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank138_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank139 (	// matmul/matmul-hw.mlir:12354:33
    .p0_rd_en   (_T_1693),	// matmul/matmul-hw.mlir:13731:13
    .p1_wr_en   (_T_1740),	// matmul/matmul-hw.mlir:13669:13
    .p1_wr_data (_T_1739),	// matmul/matmul-hw.mlir:13670:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank139_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank140 (	// matmul/matmul-hw.mlir:12355:33
    .p0_rd_en   (_T_1690),	// matmul/matmul-hw.mlir:13734:13
    .p1_wr_en   (_T_1737),	// matmul/matmul-hw.mlir:13672:13
    .p1_wr_data (_T_1736),	// matmul/matmul-hw.mlir:13673:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank140_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank141 (	// matmul/matmul-hw.mlir:12356:33
    .p0_rd_en   (_T_1687),	// matmul/matmul-hw.mlir:13737:13
    .p1_wr_en   (_T_1734),	// matmul/matmul-hw.mlir:13675:13
    .p1_wr_data (_T_1733),	// matmul/matmul-hw.mlir:13676:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank141_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank142 (	// matmul/matmul-hw.mlir:12357:33
    .p0_rd_en   (_T_1684),	// matmul/matmul-hw.mlir:13740:13
    .p1_wr_en   (_T_1731),	// matmul/matmul-hw.mlir:13678:13
    .p1_wr_data (_T_1730),	// matmul/matmul-hw.mlir:13679:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank142_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank143 (	// matmul/matmul-hw.mlir:12358:33
    .p0_rd_en   (_T_1681),	// matmul/matmul-hw.mlir:13758:13
    .p1_wr_en   (_T_1728),	// matmul/matmul-hw.mlir:13696:13
    .p1_wr_data (_T_1727),	// matmul/matmul-hw.mlir:13697:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank143_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank144 (	// matmul/matmul-hw.mlir:12359:33
    .p0_rd_en   (_T_1678),	// matmul/matmul-hw.mlir:13761:13
    .p1_wr_en   (_T_1725),	// matmul/matmul-hw.mlir:13699:13
    .p1_wr_data (_T_1724),	// matmul/matmul-hw.mlir:13700:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank144_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank145 (	// matmul/matmul-hw.mlir:12360:33
    .p0_rd_en   (_T_1675),	// matmul/matmul-hw.mlir:13764:13
    .p1_wr_en   (_T_1722),	// matmul/matmul-hw.mlir:13702:13
    .p1_wr_data (_T_1721),	// matmul/matmul-hw.mlir:13703:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank145_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank146 (	// matmul/matmul-hw.mlir:12361:33
    .p0_rd_en   (_T_1672),	// matmul/matmul-hw.mlir:13767:13
    .p1_wr_en   (_T_1719),	// matmul/matmul-hw.mlir:13705:13
    .p1_wr_data (_T_1718),	// matmul/matmul-hw.mlir:13706:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank146_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank147 (	// matmul/matmul-hw.mlir:12362:33
    .p0_rd_en   (_T_1669),	// matmul/matmul-hw.mlir:13770:13
    .p1_wr_en   (_T_1716),	// matmul/matmul-hw.mlir:13708:13
    .p1_wr_data (_T_1715),	// matmul/matmul-hw.mlir:13709:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank147_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank148 (	// matmul/matmul-hw.mlir:12363:33
    .p0_rd_en   (_T_1666),	// matmul/matmul-hw.mlir:13773:13
    .p1_wr_en   (_T_1713),	// matmul/matmul-hw.mlir:13711:13
    .p1_wr_data (_T_1712),	// matmul/matmul-hw.mlir:13712:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank148_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank149 (	// matmul/matmul-hw.mlir:12364:33
    .p0_rd_en   (_T_1663),	// matmul/matmul-hw.mlir:13776:13
    .p1_wr_en   (_T_1710),	// matmul/matmul-hw.mlir:13714:13
    .p1_wr_data (_T_1709),	// matmul/matmul-hw.mlir:13715:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank149_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank150 (	// matmul/matmul-hw.mlir:12365:33
    .p0_rd_en   (_T_1660),	// matmul/matmul-hw.mlir:13779:13
    .p1_wr_en   (_T_1707),	// matmul/matmul-hw.mlir:13717:13
    .p1_wr_data (_T_1706),	// matmul/matmul-hw.mlir:13718:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank150_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank151 (	// matmul/matmul-hw.mlir:12366:33
    .p0_rd_en   (_T_1657),	// matmul/matmul-hw.mlir:13782:13
    .p1_wr_en   (_T_1704),	// matmul/matmul-hw.mlir:13720:13
    .p1_wr_data (_T_1703),	// matmul/matmul-hw.mlir:13721:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank151_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank152 (	// matmul/matmul-hw.mlir:12367:33
    .p0_rd_en   (_T_1654),	// matmul/matmul-hw.mlir:13785:13
    .p1_wr_en   (_T_1701),	// matmul/matmul-hw.mlir:13723:13
    .p1_wr_data (_T_1700),	// matmul/matmul-hw.mlir:13724:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank152_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank153 (	// matmul/matmul-hw.mlir:12368:33
    .p0_rd_en   (_T_1651),	// matmul/matmul-hw.mlir:13788:13
    .p1_wr_en   (_T_1698),	// matmul/matmul-hw.mlir:13726:13
    .p1_wr_data (_T_1697),	// matmul/matmul-hw.mlir:13727:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank153_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank154 (	// matmul/matmul-hw.mlir:12369:33
    .p0_rd_en   (_T_1648),	// matmul/matmul-hw.mlir:13791:13
    .p1_wr_en   (_T_1695),	// matmul/matmul-hw.mlir:13729:13
    .p1_wr_data (_T_1694),	// matmul/matmul-hw.mlir:13730:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank154_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank155 (	// matmul/matmul-hw.mlir:12370:33
    .p0_rd_en   (_T_1645),	// matmul/matmul-hw.mlir:13794:13
    .p1_wr_en   (_T_1692),	// matmul/matmul-hw.mlir:13732:13
    .p1_wr_data (_T_1691),	// matmul/matmul-hw.mlir:13733:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank155_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank156 (	// matmul/matmul-hw.mlir:12371:33
    .p0_rd_en   (_T_1642),	// matmul/matmul-hw.mlir:13797:13
    .p1_wr_en   (_T_1689),	// matmul/matmul-hw.mlir:13735:13
    .p1_wr_data (_T_1688),	// matmul/matmul-hw.mlir:13736:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank156_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank157 (	// matmul/matmul-hw.mlir:12372:33
    .p0_rd_en   (_T_1639),	// matmul/matmul-hw.mlir:13800:13
    .p1_wr_en   (_T_1686),	// matmul/matmul-hw.mlir:13738:13
    .p1_wr_data (_T_1685),	// matmul/matmul-hw.mlir:13739:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank157_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank158 (	// matmul/matmul-hw.mlir:12373:33
    .p0_rd_en   (_T_1636),	// matmul/matmul-hw.mlir:13803:13
    .p1_wr_en   (_T_1683),	// matmul/matmul-hw.mlir:13741:13
    .p1_wr_data (_T_1682),	// matmul/matmul-hw.mlir:13742:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank158_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank159 (	// matmul/matmul-hw.mlir:12374:33
    .p0_rd_en   (_T_1633),	// matmul/matmul-hw.mlir:13821:13
    .p1_wr_en   (_T_1680),	// matmul/matmul-hw.mlir:13759:13
    .p1_wr_data (_T_1679),	// matmul/matmul-hw.mlir:13760:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank159_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank160 (	// matmul/matmul-hw.mlir:12375:33
    .p0_rd_en   (_T_1630),	// matmul/matmul-hw.mlir:13824:13
    .p1_wr_en   (_T_1677),	// matmul/matmul-hw.mlir:13762:13
    .p1_wr_data (_T_1676),	// matmul/matmul-hw.mlir:13763:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank160_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank161 (	// matmul/matmul-hw.mlir:12376:33
    .p0_rd_en   (_T_1627),	// matmul/matmul-hw.mlir:13827:13
    .p1_wr_en   (_T_1674),	// matmul/matmul-hw.mlir:13765:13
    .p1_wr_data (_T_1673),	// matmul/matmul-hw.mlir:13766:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank161_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank162 (	// matmul/matmul-hw.mlir:12377:33
    .p0_rd_en   (_T_1624),	// matmul/matmul-hw.mlir:13830:13
    .p1_wr_en   (_T_1671),	// matmul/matmul-hw.mlir:13768:13
    .p1_wr_data (_T_1670),	// matmul/matmul-hw.mlir:13769:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank162_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank163 (	// matmul/matmul-hw.mlir:12378:33
    .p0_rd_en   (_T_1621),	// matmul/matmul-hw.mlir:13833:13
    .p1_wr_en   (_T_1668),	// matmul/matmul-hw.mlir:13771:13
    .p1_wr_data (_T_1667),	// matmul/matmul-hw.mlir:13772:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank163_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank164 (	// matmul/matmul-hw.mlir:12379:33
    .p0_rd_en   (_T_1618),	// matmul/matmul-hw.mlir:13836:13
    .p1_wr_en   (_T_1665),	// matmul/matmul-hw.mlir:13774:13
    .p1_wr_data (_T_1664),	// matmul/matmul-hw.mlir:13775:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank164_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank165 (	// matmul/matmul-hw.mlir:12380:33
    .p0_rd_en   (_T_1615),	// matmul/matmul-hw.mlir:13839:13
    .p1_wr_en   (_T_1662),	// matmul/matmul-hw.mlir:13777:13
    .p1_wr_data (_T_1661),	// matmul/matmul-hw.mlir:13778:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank165_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank166 (	// matmul/matmul-hw.mlir:12381:33
    .p0_rd_en   (_T_1612),	// matmul/matmul-hw.mlir:13842:13
    .p1_wr_en   (_T_1659),	// matmul/matmul-hw.mlir:13780:13
    .p1_wr_data (_T_1658),	// matmul/matmul-hw.mlir:13781:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank166_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank167 (	// matmul/matmul-hw.mlir:12382:33
    .p0_rd_en   (_T_1609),	// matmul/matmul-hw.mlir:13845:13
    .p1_wr_en   (_T_1656),	// matmul/matmul-hw.mlir:13783:13
    .p1_wr_data (_T_1655),	// matmul/matmul-hw.mlir:13784:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank167_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank168 (	// matmul/matmul-hw.mlir:12383:33
    .p0_rd_en   (_T_1606),	// matmul/matmul-hw.mlir:13848:13
    .p1_wr_en   (_T_1653),	// matmul/matmul-hw.mlir:13786:13
    .p1_wr_data (_T_1652),	// matmul/matmul-hw.mlir:13787:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank168_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank169 (	// matmul/matmul-hw.mlir:12384:33
    .p0_rd_en   (_T_1603),	// matmul/matmul-hw.mlir:13851:13
    .p1_wr_en   (_T_1650),	// matmul/matmul-hw.mlir:13789:13
    .p1_wr_data (_T_1649),	// matmul/matmul-hw.mlir:13790:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank169_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank170 (	// matmul/matmul-hw.mlir:12385:33
    .p0_rd_en   (_T_1600),	// matmul/matmul-hw.mlir:13854:13
    .p1_wr_en   (_T_1647),	// matmul/matmul-hw.mlir:13792:13
    .p1_wr_data (_T_1646),	// matmul/matmul-hw.mlir:13793:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank170_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank171 (	// matmul/matmul-hw.mlir:12386:33
    .p0_rd_en   (_T_1597),	// matmul/matmul-hw.mlir:13857:13
    .p1_wr_en   (_T_1644),	// matmul/matmul-hw.mlir:13795:13
    .p1_wr_data (_T_1643),	// matmul/matmul-hw.mlir:13796:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank171_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank172 (	// matmul/matmul-hw.mlir:12387:33
    .p0_rd_en   (_T_1594),	// matmul/matmul-hw.mlir:13860:13
    .p1_wr_en   (_T_1641),	// matmul/matmul-hw.mlir:13798:13
    .p1_wr_data (_T_1640),	// matmul/matmul-hw.mlir:13799:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank172_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank173 (	// matmul/matmul-hw.mlir:12388:33
    .p0_rd_en   (_T_1591),	// matmul/matmul-hw.mlir:13863:13
    .p1_wr_en   (_T_1638),	// matmul/matmul-hw.mlir:13801:13
    .p1_wr_data (_T_1637),	// matmul/matmul-hw.mlir:13802:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank173_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank174 (	// matmul/matmul-hw.mlir:12389:33
    .p0_rd_en   (_T_1588),	// matmul/matmul-hw.mlir:13866:13
    .p1_wr_en   (_T_1635),	// matmul/matmul-hw.mlir:13804:13
    .p1_wr_data (_T_1634),	// matmul/matmul-hw.mlir:13805:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank174_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank175 (	// matmul/matmul-hw.mlir:12390:33
    .p0_rd_en   (_T_1585),	// matmul/matmul-hw.mlir:13884:13
    .p1_wr_en   (_T_1632),	// matmul/matmul-hw.mlir:13822:13
    .p1_wr_data (_T_1631),	// matmul/matmul-hw.mlir:13823:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank175_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank176 (	// matmul/matmul-hw.mlir:12391:33
    .p0_rd_en   (_T_1582),	// matmul/matmul-hw.mlir:13887:13
    .p1_wr_en   (_T_1629),	// matmul/matmul-hw.mlir:13825:13
    .p1_wr_data (_T_1628),	// matmul/matmul-hw.mlir:13826:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank176_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank177 (	// matmul/matmul-hw.mlir:12392:33
    .p0_rd_en   (_T_1579),	// matmul/matmul-hw.mlir:13890:13
    .p1_wr_en   (_T_1626),	// matmul/matmul-hw.mlir:13828:13
    .p1_wr_data (_T_1625),	// matmul/matmul-hw.mlir:13829:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank177_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank178 (	// matmul/matmul-hw.mlir:12393:33
    .p0_rd_en   (_T_1576),	// matmul/matmul-hw.mlir:13893:13
    .p1_wr_en   (_T_1623),	// matmul/matmul-hw.mlir:13831:13
    .p1_wr_data (_T_1622),	// matmul/matmul-hw.mlir:13832:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank178_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank179 (	// matmul/matmul-hw.mlir:12394:33
    .p0_rd_en   (_T_1573),	// matmul/matmul-hw.mlir:13896:13
    .p1_wr_en   (_T_1620),	// matmul/matmul-hw.mlir:13834:13
    .p1_wr_data (_T_1619),	// matmul/matmul-hw.mlir:13835:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank179_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank180 (	// matmul/matmul-hw.mlir:12395:33
    .p0_rd_en   (_T_1570),	// matmul/matmul-hw.mlir:13899:13
    .p1_wr_en   (_T_1617),	// matmul/matmul-hw.mlir:13837:13
    .p1_wr_data (_T_1616),	// matmul/matmul-hw.mlir:13838:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank180_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank181 (	// matmul/matmul-hw.mlir:12396:33
    .p0_rd_en   (_T_1567),	// matmul/matmul-hw.mlir:13902:13
    .p1_wr_en   (_T_1614),	// matmul/matmul-hw.mlir:13840:13
    .p1_wr_data (_T_1613),	// matmul/matmul-hw.mlir:13841:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank181_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank182 (	// matmul/matmul-hw.mlir:12397:33
    .p0_rd_en   (_T_1564),	// matmul/matmul-hw.mlir:13905:13
    .p1_wr_en   (_T_1611),	// matmul/matmul-hw.mlir:13843:13
    .p1_wr_data (_T_1610),	// matmul/matmul-hw.mlir:13844:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank182_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank183 (	// matmul/matmul-hw.mlir:12398:33
    .p0_rd_en   (_T_1561),	// matmul/matmul-hw.mlir:13908:13
    .p1_wr_en   (_T_1608),	// matmul/matmul-hw.mlir:13846:13
    .p1_wr_data (_T_1607),	// matmul/matmul-hw.mlir:13847:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank183_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank184 (	// matmul/matmul-hw.mlir:12399:33
    .p0_rd_en   (_T_1558),	// matmul/matmul-hw.mlir:13911:13
    .p1_wr_en   (_T_1605),	// matmul/matmul-hw.mlir:13849:13
    .p1_wr_data (_T_1604),	// matmul/matmul-hw.mlir:13850:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank184_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank185 (	// matmul/matmul-hw.mlir:12400:33
    .p0_rd_en   (_T_1555),	// matmul/matmul-hw.mlir:13914:13
    .p1_wr_en   (_T_1602),	// matmul/matmul-hw.mlir:13852:13
    .p1_wr_data (_T_1601),	// matmul/matmul-hw.mlir:13853:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank185_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank186 (	// matmul/matmul-hw.mlir:12401:33
    .p0_rd_en   (_T_1552),	// matmul/matmul-hw.mlir:13917:13
    .p1_wr_en   (_T_1599),	// matmul/matmul-hw.mlir:13855:13
    .p1_wr_data (_T_1598),	// matmul/matmul-hw.mlir:13856:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank186_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank187 (	// matmul/matmul-hw.mlir:12402:33
    .p0_rd_en   (_T_1549),	// matmul/matmul-hw.mlir:13920:13
    .p1_wr_en   (_T_1596),	// matmul/matmul-hw.mlir:13858:13
    .p1_wr_data (_T_1595),	// matmul/matmul-hw.mlir:13859:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank187_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank188 (	// matmul/matmul-hw.mlir:12403:33
    .p0_rd_en   (_T_1546),	// matmul/matmul-hw.mlir:13923:13
    .p1_wr_en   (_T_1593),	// matmul/matmul-hw.mlir:13861:13
    .p1_wr_data (_T_1592),	// matmul/matmul-hw.mlir:13862:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank188_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank189 (	// matmul/matmul-hw.mlir:12404:33
    .p0_rd_en   (_T_1543),	// matmul/matmul-hw.mlir:13926:13
    .p1_wr_en   (_T_1590),	// matmul/matmul-hw.mlir:13864:13
    .p1_wr_data (_T_1589),	// matmul/matmul-hw.mlir:13865:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank189_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank190 (	// matmul/matmul-hw.mlir:12405:33
    .p0_rd_en   (_T_1540),	// matmul/matmul-hw.mlir:13929:13
    .p1_wr_en   (_T_1587),	// matmul/matmul-hw.mlir:13867:13
    .p1_wr_data (_T_1586),	// matmul/matmul-hw.mlir:13868:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank190_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank191 (	// matmul/matmul-hw.mlir:12406:33
    .p0_rd_en   (_T_1537),	// matmul/matmul-hw.mlir:13947:13
    .p1_wr_en   (_T_1584),	// matmul/matmul-hw.mlir:13885:13
    .p1_wr_data (_T_1583),	// matmul/matmul-hw.mlir:13886:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank191_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank192 (	// matmul/matmul-hw.mlir:12407:33
    .p0_rd_en   (_T_1534),	// matmul/matmul-hw.mlir:13950:13
    .p1_wr_en   (_T_1581),	// matmul/matmul-hw.mlir:13888:13
    .p1_wr_data (_T_1580),	// matmul/matmul-hw.mlir:13889:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank192_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank193 (	// matmul/matmul-hw.mlir:12408:33
    .p0_rd_en   (_T_1531),	// matmul/matmul-hw.mlir:13953:13
    .p1_wr_en   (_T_1578),	// matmul/matmul-hw.mlir:13891:13
    .p1_wr_data (_T_1577),	// matmul/matmul-hw.mlir:13892:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank193_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank194 (	// matmul/matmul-hw.mlir:12409:33
    .p0_rd_en   (_T_1528),	// matmul/matmul-hw.mlir:13956:13
    .p1_wr_en   (_T_1575),	// matmul/matmul-hw.mlir:13894:13
    .p1_wr_data (_T_1574),	// matmul/matmul-hw.mlir:13895:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank194_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank195 (	// matmul/matmul-hw.mlir:12410:33
    .p0_rd_en   (_T_1525),	// matmul/matmul-hw.mlir:13959:13
    .p1_wr_en   (_T_1572),	// matmul/matmul-hw.mlir:13897:13
    .p1_wr_data (_T_1571),	// matmul/matmul-hw.mlir:13898:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank195_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank196 (	// matmul/matmul-hw.mlir:12411:33
    .p0_rd_en   (_T_1522),	// matmul/matmul-hw.mlir:13962:13
    .p1_wr_en   (_T_1569),	// matmul/matmul-hw.mlir:13900:13
    .p1_wr_data (_T_1568),	// matmul/matmul-hw.mlir:13901:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank196_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank197 (	// matmul/matmul-hw.mlir:12412:33
    .p0_rd_en   (_T_1519),	// matmul/matmul-hw.mlir:13965:13
    .p1_wr_en   (_T_1566),	// matmul/matmul-hw.mlir:13903:13
    .p1_wr_data (_T_1565),	// matmul/matmul-hw.mlir:13904:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank197_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank198 (	// matmul/matmul-hw.mlir:12413:33
    .p0_rd_en   (_T_1516),	// matmul/matmul-hw.mlir:13968:13
    .p1_wr_en   (_T_1563),	// matmul/matmul-hw.mlir:13906:13
    .p1_wr_data (_T_1562),	// matmul/matmul-hw.mlir:13907:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank198_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank199 (	// matmul/matmul-hw.mlir:12414:33
    .p0_rd_en   (_T_1513),	// matmul/matmul-hw.mlir:13971:13
    .p1_wr_en   (_T_1560),	// matmul/matmul-hw.mlir:13909:13
    .p1_wr_data (_T_1559),	// matmul/matmul-hw.mlir:13910:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank199_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank200 (	// matmul/matmul-hw.mlir:12415:33
    .p0_rd_en   (_T_1510),	// matmul/matmul-hw.mlir:13974:13
    .p1_wr_en   (_T_1557),	// matmul/matmul-hw.mlir:13912:13
    .p1_wr_data (_T_1556),	// matmul/matmul-hw.mlir:13913:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank200_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank201 (	// matmul/matmul-hw.mlir:12416:33
    .p0_rd_en   (_T_1507),	// matmul/matmul-hw.mlir:13977:13
    .p1_wr_en   (_T_1554),	// matmul/matmul-hw.mlir:13915:13
    .p1_wr_data (_T_1553),	// matmul/matmul-hw.mlir:13916:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank201_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank202 (	// matmul/matmul-hw.mlir:12417:33
    .p0_rd_en   (_T_1504),	// matmul/matmul-hw.mlir:13980:13
    .p1_wr_en   (_T_1551),	// matmul/matmul-hw.mlir:13918:13
    .p1_wr_data (_T_1550),	// matmul/matmul-hw.mlir:13919:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank202_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank203 (	// matmul/matmul-hw.mlir:12418:33
    .p0_rd_en   (_T_1501),	// matmul/matmul-hw.mlir:13983:13
    .p1_wr_en   (_T_1548),	// matmul/matmul-hw.mlir:13921:13
    .p1_wr_data (_T_1547),	// matmul/matmul-hw.mlir:13922:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank203_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank204 (	// matmul/matmul-hw.mlir:12419:33
    .p0_rd_en   (_T_1498),	// matmul/matmul-hw.mlir:13986:13
    .p1_wr_en   (_T_1545),	// matmul/matmul-hw.mlir:13924:13
    .p1_wr_data (_T_1544),	// matmul/matmul-hw.mlir:13925:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank204_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank205 (	// matmul/matmul-hw.mlir:12420:33
    .p0_rd_en   (_T_1495),	// matmul/matmul-hw.mlir:13989:13
    .p1_wr_en   (_T_1542),	// matmul/matmul-hw.mlir:13927:13
    .p1_wr_data (_T_1541),	// matmul/matmul-hw.mlir:13928:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank205_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank206 (	// matmul/matmul-hw.mlir:12421:33
    .p0_rd_en   (_T_1492),	// matmul/matmul-hw.mlir:13992:13
    .p1_wr_en   (_T_1539),	// matmul/matmul-hw.mlir:13930:13
    .p1_wr_data (_T_1538),	// matmul/matmul-hw.mlir:13931:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank206_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank207 (	// matmul/matmul-hw.mlir:12422:33
    .p0_rd_en   (_T_1489),	// matmul/matmul-hw.mlir:14010:13
    .p1_wr_en   (_T_1536),	// matmul/matmul-hw.mlir:13948:13
    .p1_wr_data (_T_1535),	// matmul/matmul-hw.mlir:13949:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank207_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank208 (	// matmul/matmul-hw.mlir:12423:33
    .p0_rd_en   (_T_1486),	// matmul/matmul-hw.mlir:14013:13
    .p1_wr_en   (_T_1533),	// matmul/matmul-hw.mlir:13951:13
    .p1_wr_data (_T_1532),	// matmul/matmul-hw.mlir:13952:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank208_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank209 (	// matmul/matmul-hw.mlir:12424:33
    .p0_rd_en   (_T_1483),	// matmul/matmul-hw.mlir:14016:13
    .p1_wr_en   (_T_1530),	// matmul/matmul-hw.mlir:13954:13
    .p1_wr_data (_T_1529),	// matmul/matmul-hw.mlir:13955:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank209_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank210 (	// matmul/matmul-hw.mlir:12425:33
    .p0_rd_en   (_T_1480),	// matmul/matmul-hw.mlir:14019:13
    .p1_wr_en   (_T_1527),	// matmul/matmul-hw.mlir:13957:13
    .p1_wr_data (_T_1526),	// matmul/matmul-hw.mlir:13958:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank210_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank211 (	// matmul/matmul-hw.mlir:12426:33
    .p0_rd_en   (_T_1477),	// matmul/matmul-hw.mlir:14022:13
    .p1_wr_en   (_T_1524),	// matmul/matmul-hw.mlir:13960:13
    .p1_wr_data (_T_1523),	// matmul/matmul-hw.mlir:13961:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank211_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank212 (	// matmul/matmul-hw.mlir:12427:33
    .p0_rd_en   (_T_1474),	// matmul/matmul-hw.mlir:14025:13
    .p1_wr_en   (_T_1521),	// matmul/matmul-hw.mlir:13963:13
    .p1_wr_data (_T_1520),	// matmul/matmul-hw.mlir:13964:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank212_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank213 (	// matmul/matmul-hw.mlir:12428:33
    .p0_rd_en   (_T_1471),	// matmul/matmul-hw.mlir:14028:13
    .p1_wr_en   (_T_1518),	// matmul/matmul-hw.mlir:13966:13
    .p1_wr_data (_T_1517),	// matmul/matmul-hw.mlir:13967:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank213_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank214 (	// matmul/matmul-hw.mlir:12429:33
    .p0_rd_en   (_T_1468),	// matmul/matmul-hw.mlir:14031:13
    .p1_wr_en   (_T_1515),	// matmul/matmul-hw.mlir:13969:13
    .p1_wr_data (_T_1514),	// matmul/matmul-hw.mlir:13970:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank214_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank215 (	// matmul/matmul-hw.mlir:12430:33
    .p0_rd_en   (_T_1465),	// matmul/matmul-hw.mlir:14034:13
    .p1_wr_en   (_T_1512),	// matmul/matmul-hw.mlir:13972:13
    .p1_wr_data (_T_1511),	// matmul/matmul-hw.mlir:13973:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank215_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank216 (	// matmul/matmul-hw.mlir:12431:33
    .p0_rd_en   (_T_1462),	// matmul/matmul-hw.mlir:14037:13
    .p1_wr_en   (_T_1509),	// matmul/matmul-hw.mlir:13975:13
    .p1_wr_data (_T_1508),	// matmul/matmul-hw.mlir:13976:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank216_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank217 (	// matmul/matmul-hw.mlir:12432:33
    .p0_rd_en   (_T_1459),	// matmul/matmul-hw.mlir:14040:13
    .p1_wr_en   (_T_1506),	// matmul/matmul-hw.mlir:13978:13
    .p1_wr_data (_T_1505),	// matmul/matmul-hw.mlir:13979:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank217_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank218 (	// matmul/matmul-hw.mlir:12433:33
    .p0_rd_en   (_T_1456),	// matmul/matmul-hw.mlir:14043:13
    .p1_wr_en   (_T_1503),	// matmul/matmul-hw.mlir:13981:13
    .p1_wr_data (_T_1502),	// matmul/matmul-hw.mlir:13982:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank218_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank219 (	// matmul/matmul-hw.mlir:12434:33
    .p0_rd_en   (_T_1453),	// matmul/matmul-hw.mlir:14046:13
    .p1_wr_en   (_T_1500),	// matmul/matmul-hw.mlir:13984:13
    .p1_wr_data (_T_1499),	// matmul/matmul-hw.mlir:13985:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank219_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank220 (	// matmul/matmul-hw.mlir:12435:33
    .p0_rd_en   (_T_1450),	// matmul/matmul-hw.mlir:14049:13
    .p1_wr_en   (_T_1497),	// matmul/matmul-hw.mlir:13987:13
    .p1_wr_data (_T_1496),	// matmul/matmul-hw.mlir:13988:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank220_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank221 (	// matmul/matmul-hw.mlir:12436:33
    .p0_rd_en   (_T_1447),	// matmul/matmul-hw.mlir:14052:13
    .p1_wr_en   (_T_1494),	// matmul/matmul-hw.mlir:13990:13
    .p1_wr_data (_T_1493),	// matmul/matmul-hw.mlir:13991:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank221_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank222 (	// matmul/matmul-hw.mlir:12437:33
    .p0_rd_en   (_T_1444),	// matmul/matmul-hw.mlir:14055:13
    .p1_wr_en   (_T_1491),	// matmul/matmul-hw.mlir:13993:13
    .p1_wr_data (_T_1490),	// matmul/matmul-hw.mlir:13994:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank222_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank223 (	// matmul/matmul-hw.mlir:12438:33
    .p0_rd_en   (_T_1441),	// matmul/matmul-hw.mlir:14073:13
    .p1_wr_en   (_T_1488),	// matmul/matmul-hw.mlir:14011:13
    .p1_wr_data (_T_1487),	// matmul/matmul-hw.mlir:14012:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank223_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank224 (	// matmul/matmul-hw.mlir:12439:33
    .p0_rd_en   (_T_1438),	// matmul/matmul-hw.mlir:14076:13
    .p1_wr_en   (_T_1485),	// matmul/matmul-hw.mlir:14014:13
    .p1_wr_data (_T_1484),	// matmul/matmul-hw.mlir:14015:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank224_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank225 (	// matmul/matmul-hw.mlir:12440:33
    .p0_rd_en   (_T_1435),	// matmul/matmul-hw.mlir:14079:13
    .p1_wr_en   (_T_1482),	// matmul/matmul-hw.mlir:14017:13
    .p1_wr_data (_T_1481),	// matmul/matmul-hw.mlir:14018:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank225_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank226 (	// matmul/matmul-hw.mlir:12441:33
    .p0_rd_en   (_T_1432),	// matmul/matmul-hw.mlir:14082:13
    .p1_wr_en   (_T_1479),	// matmul/matmul-hw.mlir:14020:13
    .p1_wr_data (_T_1478),	// matmul/matmul-hw.mlir:14021:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank226_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank227 (	// matmul/matmul-hw.mlir:12442:33
    .p0_rd_en   (_T_1429),	// matmul/matmul-hw.mlir:14085:13
    .p1_wr_en   (_T_1476),	// matmul/matmul-hw.mlir:14023:13
    .p1_wr_data (_T_1475),	// matmul/matmul-hw.mlir:14024:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank227_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank228 (	// matmul/matmul-hw.mlir:12443:33
    .p0_rd_en   (_T_1426),	// matmul/matmul-hw.mlir:14088:13
    .p1_wr_en   (_T_1473),	// matmul/matmul-hw.mlir:14026:13
    .p1_wr_data (_T_1472),	// matmul/matmul-hw.mlir:14027:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank228_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank229 (	// matmul/matmul-hw.mlir:12444:33
    .p0_rd_en   (_T_1423),	// matmul/matmul-hw.mlir:14091:13
    .p1_wr_en   (_T_1470),	// matmul/matmul-hw.mlir:14029:13
    .p1_wr_data (_T_1469),	// matmul/matmul-hw.mlir:14030:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank229_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank230 (	// matmul/matmul-hw.mlir:12445:33
    .p0_rd_en   (_T_1420),	// matmul/matmul-hw.mlir:14094:13
    .p1_wr_en   (_T_1467),	// matmul/matmul-hw.mlir:14032:13
    .p1_wr_data (_T_1466),	// matmul/matmul-hw.mlir:14033:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank230_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank231 (	// matmul/matmul-hw.mlir:12446:33
    .p0_rd_en   (_T_1417),	// matmul/matmul-hw.mlir:14097:13
    .p1_wr_en   (_T_1464),	// matmul/matmul-hw.mlir:14035:13
    .p1_wr_data (_T_1463),	// matmul/matmul-hw.mlir:14036:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank231_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank232 (	// matmul/matmul-hw.mlir:12447:33
    .p0_rd_en   (_T_1414),	// matmul/matmul-hw.mlir:14100:13
    .p1_wr_en   (_T_1461),	// matmul/matmul-hw.mlir:14038:13
    .p1_wr_data (_T_1460),	// matmul/matmul-hw.mlir:14039:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank232_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank233 (	// matmul/matmul-hw.mlir:12448:33
    .p0_rd_en   (_T_1411),	// matmul/matmul-hw.mlir:14103:13
    .p1_wr_en   (_T_1458),	// matmul/matmul-hw.mlir:14041:13
    .p1_wr_data (_T_1457),	// matmul/matmul-hw.mlir:14042:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank233_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank234 (	// matmul/matmul-hw.mlir:12449:33
    .p0_rd_en   (_T_1408),	// matmul/matmul-hw.mlir:14106:13
    .p1_wr_en   (_T_1455),	// matmul/matmul-hw.mlir:14044:13
    .p1_wr_data (_T_1454),	// matmul/matmul-hw.mlir:14045:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank234_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank235 (	// matmul/matmul-hw.mlir:12450:33
    .p0_rd_en   (_T_1405),	// matmul/matmul-hw.mlir:14109:13
    .p1_wr_en   (_T_1452),	// matmul/matmul-hw.mlir:14047:13
    .p1_wr_data (_T_1451),	// matmul/matmul-hw.mlir:14048:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank235_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank236 (	// matmul/matmul-hw.mlir:12451:33
    .p0_rd_en   (_T_1402),	// matmul/matmul-hw.mlir:14112:13
    .p1_wr_en   (_T_1449),	// matmul/matmul-hw.mlir:14050:13
    .p1_wr_data (_T_1448),	// matmul/matmul-hw.mlir:14051:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank236_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank237 (	// matmul/matmul-hw.mlir:12452:33
    .p0_rd_en   (_T_1399),	// matmul/matmul-hw.mlir:14115:13
    .p1_wr_en   (_T_1446),	// matmul/matmul-hw.mlir:14053:13
    .p1_wr_data (_T_1445),	// matmul/matmul-hw.mlir:14054:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank237_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank238 (	// matmul/matmul-hw.mlir:12453:33
    .p0_rd_en   (_T_1396),	// matmul/matmul-hw.mlir:14118:13
    .p1_wr_en   (_T_1443),	// matmul/matmul-hw.mlir:14056:13
    .p1_wr_data (_T_1442),	// matmul/matmul-hw.mlir:14057:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank238_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank239 (	// matmul/matmul-hw.mlir:12454:33
    .p0_rd_en   (_T_1393),	// matmul/matmul-hw.mlir:14136:13
    .p1_wr_en   (_T_1440),	// matmul/matmul-hw.mlir:14074:13
    .p1_wr_data (_T_1439),	// matmul/matmul-hw.mlir:14075:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank239_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank240 (	// matmul/matmul-hw.mlir:12455:33
    .p0_rd_en   (_T_83),	// matmul/matmul-hw.mlir:23068:13
    .p1_wr_en   (_T_1437),	// matmul/matmul-hw.mlir:14077:13
    .p1_wr_data (_T_1436),	// matmul/matmul-hw.mlir:14078:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank240_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank241 (	// matmul/matmul-hw.mlir:12456:33
    .p0_rd_en   (_T_78),	// matmul/matmul-hw.mlir:23098:13
    .p1_wr_en   (_T_1434),	// matmul/matmul-hw.mlir:14080:13
    .p1_wr_data (_T_1433),	// matmul/matmul-hw.mlir:14081:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank241_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank242 (	// matmul/matmul-hw.mlir:12457:33
    .p0_rd_en   (_T_73),	// matmul/matmul-hw.mlir:23128:13
    .p1_wr_en   (_T_1431),	// matmul/matmul-hw.mlir:14083:13
    .p1_wr_data (_T_1430),	// matmul/matmul-hw.mlir:14084:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank242_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank243 (	// matmul/matmul-hw.mlir:12458:33
    .p0_rd_en   (_T_68),	// matmul/matmul-hw.mlir:23158:13
    .p1_wr_en   (_T_1428),	// matmul/matmul-hw.mlir:14086:13
    .p1_wr_data (_T_1427),	// matmul/matmul-hw.mlir:14087:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank243_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank244 (	// matmul/matmul-hw.mlir:12459:33
    .p0_rd_en   (_T_63),	// matmul/matmul-hw.mlir:23188:13
    .p1_wr_en   (_T_1425),	// matmul/matmul-hw.mlir:14089:13
    .p1_wr_data (_T_1424),	// matmul/matmul-hw.mlir:14090:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank244_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank245 (	// matmul/matmul-hw.mlir:12460:33
    .p0_rd_en   (_T_58),	// matmul/matmul-hw.mlir:23218:13
    .p1_wr_en   (_T_1422),	// matmul/matmul-hw.mlir:14092:13
    .p1_wr_data (_T_1421),	// matmul/matmul-hw.mlir:14093:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank245_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank246 (	// matmul/matmul-hw.mlir:12461:33
    .p0_rd_en   (_T_53),	// matmul/matmul-hw.mlir:23248:13
    .p1_wr_en   (_T_1419),	// matmul/matmul-hw.mlir:14095:13
    .p1_wr_data (_T_1418),	// matmul/matmul-hw.mlir:14096:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank246_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank247 (	// matmul/matmul-hw.mlir:12462:33
    .p0_rd_en   (_T_48),	// matmul/matmul-hw.mlir:23278:13
    .p1_wr_en   (_T_1416),	// matmul/matmul-hw.mlir:14098:13
    .p1_wr_data (_T_1415),	// matmul/matmul-hw.mlir:14099:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank247_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank248 (	// matmul/matmul-hw.mlir:12463:33
    .p0_rd_en   (_T_43),	// matmul/matmul-hw.mlir:23308:13
    .p1_wr_en   (_T_1413),	// matmul/matmul-hw.mlir:14101:13
    .p1_wr_data (_T_1412),	// matmul/matmul-hw.mlir:14102:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank248_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank249 (	// matmul/matmul-hw.mlir:12464:33
    .p0_rd_en   (_T_38),	// matmul/matmul-hw.mlir:23338:13
    .p1_wr_en   (_T_1410),	// matmul/matmul-hw.mlir:14104:13
    .p1_wr_data (_T_1409),	// matmul/matmul-hw.mlir:14105:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank249_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank250 (	// matmul/matmul-hw.mlir:12465:33
    .p0_rd_en   (_T_33),	// matmul/matmul-hw.mlir:23368:13
    .p1_wr_en   (_T_1407),	// matmul/matmul-hw.mlir:14107:13
    .p1_wr_data (_T_1406),	// matmul/matmul-hw.mlir:14108:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank250_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank251 (	// matmul/matmul-hw.mlir:12466:33
    .p0_rd_en   (_T_28),	// matmul/matmul-hw.mlir:23398:13
    .p1_wr_en   (_T_1404),	// matmul/matmul-hw.mlir:14110:13
    .p1_wr_data (_T_1403),	// matmul/matmul-hw.mlir:14111:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank251_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank252 (	// matmul/matmul-hw.mlir:12467:33
    .p0_rd_en   (_T_23),	// matmul/matmul-hw.mlir:23428:13
    .p1_wr_en   (_T_1401),	// matmul/matmul-hw.mlir:14113:13
    .p1_wr_data (_T_1400),	// matmul/matmul-hw.mlir:14114:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank252_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank253 (	// matmul/matmul-hw.mlir:12468:33
    .p0_rd_en   (_T_18),	// matmul/matmul-hw.mlir:23458:13
    .p1_wr_en   (_T_1398),	// matmul/matmul-hw.mlir:14116:13
    .p1_wr_data (_T_1397),	// matmul/matmul-hw.mlir:14117:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank253_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank254 (	// matmul/matmul-hw.mlir:12469:33
    .p0_rd_en   (_T_13),	// matmul/matmul-hw.mlir:23488:13
    .p1_wr_en   (_T_1395),	// matmul/matmul-hw.mlir:14119:13
    .p1_wr_data (_T_1394),	// matmul/matmul-hw.mlir:14120:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank254_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) A_reg_bank255 (	// matmul/matmul-hw.mlir:12470:33
    .p0_rd_en   (_T_8),	// matmul/matmul-hw.mlir:23518:13
    .p1_wr_en   (_T_1392),	// matmul/matmul-hw.mlir:14137:13
    .p1_wr_data (_T_1391),	// matmul/matmul-hw.mlir:14138:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (A_reg_bank255_p0_rd_data)
  );
  wire [3:0] _T_2718 = _T_2717[3:0];	// matmul/matmul-hw.mlir:12471:12
  assign _T_2192 = _T_2712 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12472:12
  assign _T_2191 = _T_2712 ? _T_2718 : 4'bx;	// matmul/matmul-hw.mlir:10224:18, :12473:12
  assign _T_2190 = _T_2712 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12474:12
  localparam _T_2720 = 1'h0;	// matmul/matmul-hw.mlir:12477:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12478:5
    if (rst)	// matmul/matmul-hw.mlir:12478:5
      _T_2719 <= _T_2720;	// matmul/matmul-hw.mlir:12481:7
    else	// matmul/matmul-hw.mlir:12478:5
      _T_2719 <= _T_2712;	// matmul/matmul-hw.mlir:12479:7
  end // always @(posedge)
  assign _T_2188 = _T_2189;	// matmul/matmul-hw.mlir:12484:12
  localparam _T_2721 = 1'h0;	// matmul/matmul-hw.mlir:12485:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12486:5
    if (rst)	// matmul/matmul-hw.mlir:12486:5
      _T_2189 <= _T_2721;	// matmul/matmul-hw.mlir:12489:7
    else	// matmul/matmul-hw.mlir:12486:5
      _T_2189 <= _T_2712;	// matmul/matmul-hw.mlir:12487:7
  end // always @(posedge)
  assign _T_2187 = _T_2189 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12484:12, :12491:12
  assign _T_2186 = _T_2189 ? A_p0_rd_data[4'h0] : 32'bx;	// matmul/matmul-hw.mlir:10221:19, :11067:14, :11068:12, :12484:12, :12492:12
  localparam [3:0] _T_2722 = 4'h0;	// matmul/matmul-hw.mlir:12495:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12496:5
    if (rst)	// matmul/matmul-hw.mlir:12496:5
      i_k_next <= _T_2722;	// matmul/matmul-hw.mlir:12499:7
    else	// matmul/matmul-hw.mlir:12496:5
      i_k_next <= _T_2718;	// matmul/matmul-hw.mlir:12497:7
  end // always @(posedge)
  assign i_k_next_i_k_0 = i_k_next;	// matmul/matmul-hw.mlir:12494:12, :12502:5
  //PROBE: i_k_next_i_k_0	// matmul/matmul-hw.mlir:12503:5
  assign _T_2185 = _T_2189 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12484:12, :12504:12
  assign _T_2184 = _T_2189 ? i_k_next : 4'bx;	// matmul/matmul-hw.mlir:10219:18, :12484:12, :12494:12, :12505:12
  assign _T_2183 = _T_2189 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12484:12, :12506:12
  wire [1:0] _T_2724 = _T_2723;	// matmul/matmul-hw.mlir:12508:12
  wire [1:0] _T_2725 = {_T_2724[1'h0+:1], {{_T_2712}}};	// matmul/matmul-hw.mlir:12509:19, :12510:12, :12511:12, :12512:12
  wire [1:0] _T_2726 = {{1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12513:19, :12514:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12515:5
    if (rst)	// matmul/matmul-hw.mlir:12515:5
      _T_2723 <= _T_2726;	// matmul/matmul-hw.mlir:12518:7
    else	// matmul/matmul-hw.mlir:12515:5
      _T_2723 <= _T_2725;	// matmul/matmul-hw.mlir:12516:7
  end // always @(posedge)
  wire [1:0] _T_2728 = _T_2727;	// matmul/matmul-hw.mlir:12523:12
  wire [1:0] _T_2729 = {_T_2728[1'h0+:1], {{_T_2712}}};	// matmul/matmul-hw.mlir:12524:19, :12525:12, :12526:12, :12527:12
  wire [1:0] _T_2730 = {{1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12528:19, :12529:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12530:5
    if (rst)	// matmul/matmul-hw.mlir:12530:5
      _T_2727 <= _T_2730;	// matmul/matmul-hw.mlir:12533:7
    else	// matmul/matmul-hw.mlir:12530:5
      _T_2727 <= _T_2729;	// matmul/matmul-hw.mlir:12531:7
  end // always @(posedge)
  wire _T_2731 = _T_2727[1'h1];	// matmul/matmul-hw.mlir:12523:12, :12535:18, :12536:12
  assign _T_2182 = _T_2731 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12537:12
  assign _T_2181 = _T_2731 ? A_p0_rd_data[4'h1] : 32'bx;	// matmul/matmul-hw.mlir:10216:19, :11072:14, :11073:12, :12538:12
  localparam [3:0] _T_2733 = 4'h0;	// matmul/matmul-hw.mlir:12541:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12542:5
    if (rst)	// matmul/matmul-hw.mlir:12542:5
      i_k_next_2732 <= _T_2733;	// matmul/matmul-hw.mlir:12545:7
    else	// matmul/matmul-hw.mlir:12542:5
      i_k_next_2732 <= i_k_next;	// matmul/matmul-hw.mlir:12494:12, :12543:7
  end // always @(posedge)
  assign i_k_next_i_k_1 = i_k_next_2732;	// matmul/matmul-hw.mlir:12540:12, :12548:5
  //PROBE: i_k_next_i_k_1	// matmul/matmul-hw.mlir:12549:5
  assign _T_2180 = _T_2731 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12550:12
  assign _T_2179 = _T_2731 ? i_k_next_2732 : 4'bx;	// matmul/matmul-hw.mlir:10214:18, :12540:12, :12551:12
  assign _T_2178 = _T_2731 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12552:12
  wire [2:0] _T_2735 = _T_2734;	// matmul/matmul-hw.mlir:12554:12
  wire [2:0] _T_2736 = {_T_2735[2'h0+:2], {{_T_2712}}};	// matmul/matmul-hw.mlir:12555:14, :12556:12, :12557:12, :12558:12
  wire [2:0] _T_2737 = {{1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12559:19, :12560:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12561:5
    if (rst)	// matmul/matmul-hw.mlir:12561:5
      _T_2734 <= _T_2737;	// matmul/matmul-hw.mlir:12564:7
    else	// matmul/matmul-hw.mlir:12561:5
      _T_2734 <= _T_2736;	// matmul/matmul-hw.mlir:12562:7
  end // always @(posedge)
  wire [2:0] _T_2739 = _T_2738;	// matmul/matmul-hw.mlir:12569:12
  wire [2:0] _T_2740 = {_T_2739[2'h0+:2], {{_T_2712}}};	// matmul/matmul-hw.mlir:12570:19, :12571:12, :12572:12, :12573:12
  wire [2:0] _T_2741 = {{1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12574:19, :12575:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12576:5
    if (rst)	// matmul/matmul-hw.mlir:12576:5
      _T_2738 <= _T_2741;	// matmul/matmul-hw.mlir:12579:7
    else	// matmul/matmul-hw.mlir:12576:5
      _T_2738 <= _T_2740;	// matmul/matmul-hw.mlir:12577:7
  end // always @(posedge)
  wire _T_2742 = _T_2738[2'h2];	// matmul/matmul-hw.mlir:12569:12, :12581:20, :12582:12
  assign _T_2177 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12583:12
  assign _T_2176 = _T_2742 ? A_p0_rd_data[4'h2] : 32'bx;	// matmul/matmul-hw.mlir:10211:19, :11077:14, :11078:12, :12584:12
  localparam [3:0] _T_2744 = 4'h0;	// matmul/matmul-hw.mlir:12587:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12588:5
    if (rst)	// matmul/matmul-hw.mlir:12588:5
      i_k_next_2743 <= _T_2744;	// matmul/matmul-hw.mlir:12591:7
    else	// matmul/matmul-hw.mlir:12588:5
      i_k_next_2743 <= i_k_next_2732;	// matmul/matmul-hw.mlir:12540:12, :12589:7
  end // always @(posedge)
  assign i_k_next_i_k_2 = i_k_next_2743;	// matmul/matmul-hw.mlir:12586:12, :12594:5
  //PROBE: i_k_next_i_k_2	// matmul/matmul-hw.mlir:12595:5
  assign _T_2175 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12596:12
  assign _T_2174 = _T_2742 ? i_k_next_2743 : 4'bx;	// matmul/matmul-hw.mlir:10209:18, :12586:12, :12597:12
  assign _T_2173 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12598:12
  wire [3:0] _T_2746 = _T_2745;	// matmul/matmul-hw.mlir:12600:12
  wire [3:0] _T_2747 = {_T_2746[2'h0+:3], {{_T_2712}}};	// matmul/matmul-hw.mlir:12601:19, :12602:12, :12603:12, :12604:12
  wire [3:0] _T_2748 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12605:19, :12606:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12607:5
    if (rst)	// matmul/matmul-hw.mlir:12607:5
      _T_2745 <= _T_2748;	// matmul/matmul-hw.mlir:12610:7
    else	// matmul/matmul-hw.mlir:12607:5
      _T_2745 <= _T_2747;	// matmul/matmul-hw.mlir:12608:7
  end // always @(posedge)
  wire [3:0] _T_2750 = _T_2749;	// matmul/matmul-hw.mlir:12615:12
  wire [3:0] _T_2751 = {_T_2750[2'h0+:3], {{_T_2712}}};	// matmul/matmul-hw.mlir:12616:19, :12617:12, :12618:12, :12619:12
  wire [3:0] _T_2752 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12620:19, :12621:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12622:5
    if (rst)	// matmul/matmul-hw.mlir:12622:5
      _T_2749 <= _T_2752;	// matmul/matmul-hw.mlir:12625:7
    else	// matmul/matmul-hw.mlir:12622:5
      _T_2749 <= _T_2751;	// matmul/matmul-hw.mlir:12623:7
  end // always @(posedge)
  wire _T_2753 = _T_2749[2'h3];	// matmul/matmul-hw.mlir:12615:12, :12627:20, :12628:12
  assign _T_2172 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12629:12
  assign _T_2171 = _T_2753 ? A_p0_rd_data[4'h3] : 32'bx;	// matmul/matmul-hw.mlir:10206:19, :11082:14, :11083:12, :12630:12
  localparam [3:0] _T_2755 = 4'h0;	// matmul/matmul-hw.mlir:12633:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12634:5
    if (rst)	// matmul/matmul-hw.mlir:12634:5
      i_k_next_2754 <= _T_2755;	// matmul/matmul-hw.mlir:12637:7
    else	// matmul/matmul-hw.mlir:12634:5
      i_k_next_2754 <= i_k_next_2743;	// matmul/matmul-hw.mlir:12586:12, :12635:7
  end // always @(posedge)
  assign i_k_next_i_k_3 = i_k_next_2754;	// matmul/matmul-hw.mlir:12632:12, :12640:5
  //PROBE: i_k_next_i_k_3	// matmul/matmul-hw.mlir:12641:5
  assign _T_2170 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12642:12
  assign _T_2169 = _T_2753 ? i_k_next_2754 : 4'bx;	// matmul/matmul-hw.mlir:10204:18, :12632:12, :12643:12
  assign _T_2168 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12644:12
  wire [4:0] _T_2757 = _T_2756;	// matmul/matmul-hw.mlir:12646:12
  wire [4:0] _T_2758 = {_T_2757[3'h0+:4], {{_T_2712}}};	// matmul/matmul-hw.mlir:12647:14, :12648:12, :12649:12, :12650:12
  wire [4:0] _T_2759 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12651:19, :12652:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12653:5
    if (rst)	// matmul/matmul-hw.mlir:12653:5
      _T_2756 <= _T_2759;	// matmul/matmul-hw.mlir:12656:7
    else	// matmul/matmul-hw.mlir:12653:5
      _T_2756 <= _T_2758;	// matmul/matmul-hw.mlir:12654:7
  end // always @(posedge)
  wire [4:0] _T_2761 = _T_2760;	// matmul/matmul-hw.mlir:12661:12
  wire [4:0] _T_2762 = {_T_2761[3'h0+:4], {{_T_2712}}};	// matmul/matmul-hw.mlir:12662:19, :12663:12, :12664:12, :12665:12
  wire [4:0] _T_2763 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12666:19, :12667:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12668:5
    if (rst)	// matmul/matmul-hw.mlir:12668:5
      _T_2760 <= _T_2763;	// matmul/matmul-hw.mlir:12671:7
    else	// matmul/matmul-hw.mlir:12668:5
      _T_2760 <= _T_2762;	// matmul/matmul-hw.mlir:12669:7
  end // always @(posedge)
  wire _T_2764 = _T_2760[3'h4];	// matmul/matmul-hw.mlir:12661:12, :12673:20, :12674:12
  assign _T_2167 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12675:12
  assign _T_2166 = _T_2764 ? A_p0_rd_data[4'h4] : 32'bx;	// matmul/matmul-hw.mlir:10201:19, :11087:14, :11088:12, :12676:12
  localparam [3:0] _T_2766 = 4'h0;	// matmul/matmul-hw.mlir:12679:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12680:5
    if (rst)	// matmul/matmul-hw.mlir:12680:5
      i_k_next_2765 <= _T_2766;	// matmul/matmul-hw.mlir:12683:7
    else	// matmul/matmul-hw.mlir:12680:5
      i_k_next_2765 <= i_k_next_2754;	// matmul/matmul-hw.mlir:12632:12, :12681:7
  end // always @(posedge)
  assign i_k_next_i_k_4 = i_k_next_2765;	// matmul/matmul-hw.mlir:12678:12, :12686:5
  //PROBE: i_k_next_i_k_4	// matmul/matmul-hw.mlir:12687:5
  assign _T_2165 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12688:12
  assign _T_2164 = _T_2764 ? i_k_next_2765 : 4'bx;	// matmul/matmul-hw.mlir:10199:18, :12678:12, :12689:12
  assign _T_2163 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12690:12
  wire [5:0] _T_2768 = _T_2767;	// matmul/matmul-hw.mlir:12692:12
  wire [5:0] _T_2769 = {_T_2768[3'h0+:5], {{_T_2712}}};	// matmul/matmul-hw.mlir:12693:19, :12694:12, :12695:12, :12696:12
  wire [5:0] _T_2770 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12697:19, :12698:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12699:5
    if (rst)	// matmul/matmul-hw.mlir:12699:5
      _T_2767 <= _T_2770;	// matmul/matmul-hw.mlir:12702:7
    else	// matmul/matmul-hw.mlir:12699:5
      _T_2767 <= _T_2769;	// matmul/matmul-hw.mlir:12700:7
  end // always @(posedge)
  wire [5:0] _T_2772 = _T_2771;	// matmul/matmul-hw.mlir:12707:12
  wire [5:0] _T_2773 = {_T_2772[3'h0+:5], {{_T_2712}}};	// matmul/matmul-hw.mlir:12708:19, :12709:12, :12710:12, :12711:12
  wire [5:0] _T_2774 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12712:19, :12713:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12714:5
    if (rst)	// matmul/matmul-hw.mlir:12714:5
      _T_2771 <= _T_2774;	// matmul/matmul-hw.mlir:12717:7
    else	// matmul/matmul-hw.mlir:12714:5
      _T_2771 <= _T_2773;	// matmul/matmul-hw.mlir:12715:7
  end // always @(posedge)
  wire _T_2775 = _T_2771[3'h5];	// matmul/matmul-hw.mlir:12707:12, :12719:20, :12720:12
  assign _T_2162 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12721:12
  assign _T_2161 = _T_2775 ? A_p0_rd_data[4'h5] : 32'bx;	// matmul/matmul-hw.mlir:10196:19, :11092:14, :11093:12, :12722:12
  localparam [3:0] _T_2777 = 4'h0;	// matmul/matmul-hw.mlir:12725:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12726:5
    if (rst)	// matmul/matmul-hw.mlir:12726:5
      i_k_next_2776 <= _T_2777;	// matmul/matmul-hw.mlir:12729:7
    else	// matmul/matmul-hw.mlir:12726:5
      i_k_next_2776 <= i_k_next_2765;	// matmul/matmul-hw.mlir:12678:12, :12727:7
  end // always @(posedge)
  assign i_k_next_i_k_5 = i_k_next_2776;	// matmul/matmul-hw.mlir:12724:12, :12732:5
  //PROBE: i_k_next_i_k_5	// matmul/matmul-hw.mlir:12733:5
  assign _T_2160 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12734:12
  assign _T_2159 = _T_2775 ? i_k_next_2776 : 4'bx;	// matmul/matmul-hw.mlir:10194:18, :12724:12, :12735:12
  assign _T_2158 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12736:12
  wire [6:0] _T_2779 = _T_2778;	// matmul/matmul-hw.mlir:12738:12
  wire [6:0] _T_2780 = {_T_2779[3'h0+:6], {{_T_2712}}};	// matmul/matmul-hw.mlir:12739:19, :12740:12, :12741:12, :12742:12
  wire [6:0] _T_2781 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12743:19, :12744:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12745:5
    if (rst)	// matmul/matmul-hw.mlir:12745:5
      _T_2778 <= _T_2781;	// matmul/matmul-hw.mlir:12748:7
    else	// matmul/matmul-hw.mlir:12745:5
      _T_2778 <= _T_2780;	// matmul/matmul-hw.mlir:12746:7
  end // always @(posedge)
  wire [6:0] _T_2783 = _T_2782;	// matmul/matmul-hw.mlir:12753:12
  wire [6:0] _T_2784 = {_T_2783[3'h0+:6], {{_T_2712}}};	// matmul/matmul-hw.mlir:12754:19, :12755:12, :12756:12, :12757:12
  wire [6:0] _T_2785 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12758:19, :12759:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12760:5
    if (rst)	// matmul/matmul-hw.mlir:12760:5
      _T_2782 <= _T_2785;	// matmul/matmul-hw.mlir:12763:7
    else	// matmul/matmul-hw.mlir:12760:5
      _T_2782 <= _T_2784;	// matmul/matmul-hw.mlir:12761:7
  end // always @(posedge)
  wire _T_2786 = _T_2782[3'h6];	// matmul/matmul-hw.mlir:12753:12, :12765:20, :12766:12
  assign _T_2157 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12767:12
  assign _T_2156 = _T_2786 ? A_p0_rd_data[4'h6] : 32'bx;	// matmul/matmul-hw.mlir:10191:19, :11097:14, :11098:12, :12768:12
  localparam [3:0] _T_2788 = 4'h0;	// matmul/matmul-hw.mlir:12771:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12772:5
    if (rst)	// matmul/matmul-hw.mlir:12772:5
      i_k_next_2787 <= _T_2788;	// matmul/matmul-hw.mlir:12775:7
    else	// matmul/matmul-hw.mlir:12772:5
      i_k_next_2787 <= i_k_next_2776;	// matmul/matmul-hw.mlir:12724:12, :12773:7
  end // always @(posedge)
  assign i_k_next_i_k_6 = i_k_next_2787;	// matmul/matmul-hw.mlir:12770:12, :12778:5
  //PROBE: i_k_next_i_k_6	// matmul/matmul-hw.mlir:12779:5
  assign _T_2155 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12780:12
  assign _T_2154 = _T_2786 ? i_k_next_2787 : 4'bx;	// matmul/matmul-hw.mlir:10189:18, :12770:12, :12781:12
  assign _T_2153 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12782:12
  wire [7:0] _T_2790 = _T_2789;	// matmul/matmul-hw.mlir:12784:12
  wire [7:0] _T_2791 = {_T_2790[3'h0+:7], {{_T_2712}}};	// matmul/matmul-hw.mlir:12785:19, :12786:12, :12787:12, :12788:12
  wire [7:0] _T_2792 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12789:19, :12790:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12791:5
    if (rst)	// matmul/matmul-hw.mlir:12791:5
      _T_2789 <= _T_2792;	// matmul/matmul-hw.mlir:12794:7
    else	// matmul/matmul-hw.mlir:12791:5
      _T_2789 <= _T_2791;	// matmul/matmul-hw.mlir:12792:7
  end // always @(posedge)
  wire [7:0] _T_2794 = _T_2793;	// matmul/matmul-hw.mlir:12799:12
  wire [7:0] _T_2795 = {_T_2794[3'h0+:7], {{_T_2712}}};	// matmul/matmul-hw.mlir:12800:19, :12801:12, :12802:12, :12803:12
  wire [7:0] _T_2796 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12804:19, :12805:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12806:5
    if (rst)	// matmul/matmul-hw.mlir:12806:5
      _T_2793 <= _T_2796;	// matmul/matmul-hw.mlir:12809:7
    else	// matmul/matmul-hw.mlir:12806:5
      _T_2793 <= _T_2795;	// matmul/matmul-hw.mlir:12807:7
  end // always @(posedge)
  wire _T_2797 = _T_2793[3'h7];	// matmul/matmul-hw.mlir:12799:12, :12811:20, :12812:12
  assign _T_2152 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12813:12
  assign _T_2151 = _T_2797 ? A_p0_rd_data[4'h7] : 32'bx;	// matmul/matmul-hw.mlir:10186:19, :11102:14, :11103:12, :12814:12
  localparam [3:0] _T_2799 = 4'h0;	// matmul/matmul-hw.mlir:12817:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12818:5
    if (rst)	// matmul/matmul-hw.mlir:12818:5
      i_k_next_2798 <= _T_2799;	// matmul/matmul-hw.mlir:12821:7
    else	// matmul/matmul-hw.mlir:12818:5
      i_k_next_2798 <= i_k_next_2787;	// matmul/matmul-hw.mlir:12770:12, :12819:7
  end // always @(posedge)
  assign i_k_next_i_k_7 = i_k_next_2798;	// matmul/matmul-hw.mlir:12816:12, :12824:5
  //PROBE: i_k_next_i_k_7	// matmul/matmul-hw.mlir:12825:5
  assign _T_2150 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12826:12
  assign _T_2149 = _T_2797 ? i_k_next_2798 : 4'bx;	// matmul/matmul-hw.mlir:10184:18, :12816:12, :12827:12
  assign _T_2148 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12828:12
  wire [8:0] _T_2801 = _T_2800;	// matmul/matmul-hw.mlir:12830:12
  wire [8:0] _T_2802 = {_T_2801[4'h0+:8], {{_T_2712}}};	// matmul/matmul-hw.mlir:12831:19, :12832:12, :12833:12, :12834:12
  wire [8:0] _T_2803 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12835:19, :12836:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12837:5
    if (rst)	// matmul/matmul-hw.mlir:12837:5
      _T_2800 <= _T_2803;	// matmul/matmul-hw.mlir:12840:7
    else	// matmul/matmul-hw.mlir:12837:5
      _T_2800 <= _T_2802;	// matmul/matmul-hw.mlir:12838:7
  end // always @(posedge)
  wire [8:0] _T_2805 = _T_2804;	// matmul/matmul-hw.mlir:12845:12
  wire [8:0] _T_2806 = {_T_2805[4'h0+:8], {{_T_2712}}};	// matmul/matmul-hw.mlir:12846:19, :12847:12, :12848:12, :12849:12
  wire [8:0] _T_2807 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12850:19, :12851:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12852:5
    if (rst)	// matmul/matmul-hw.mlir:12852:5
      _T_2804 <= _T_2807;	// matmul/matmul-hw.mlir:12855:7
    else	// matmul/matmul-hw.mlir:12852:5
      _T_2804 <= _T_2806;	// matmul/matmul-hw.mlir:12853:7
  end // always @(posedge)
  wire _T_2808 = _T_2804[4'h8];	// matmul/matmul-hw.mlir:12845:12, :12857:20, :12858:12
  assign _T_2147 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12859:12
  assign _T_2146 = _T_2808 ? A_p0_rd_data[4'h8] : 32'bx;	// matmul/matmul-hw.mlir:10181:19, :11107:15, :11108:12, :12860:12
  localparam [3:0] _T_2810 = 4'h0;	// matmul/matmul-hw.mlir:12863:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12864:5
    if (rst)	// matmul/matmul-hw.mlir:12864:5
      i_k_next_2809 <= _T_2810;	// matmul/matmul-hw.mlir:12867:7
    else	// matmul/matmul-hw.mlir:12864:5
      i_k_next_2809 <= i_k_next_2798;	// matmul/matmul-hw.mlir:12816:12, :12865:7
  end // always @(posedge)
  assign i_k_next_i_k_8 = i_k_next_2809;	// matmul/matmul-hw.mlir:12862:12, :12870:5
  //PROBE: i_k_next_i_k_8	// matmul/matmul-hw.mlir:12871:5
  assign _T_2145 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12872:12
  assign _T_2144 = _T_2808 ? i_k_next_2809 : 4'bx;	// matmul/matmul-hw.mlir:10179:18, :12862:12, :12873:12
  assign _T_2143 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12874:12
  wire [9:0] _T_2812 = _T_2811;	// matmul/matmul-hw.mlir:12876:12
  wire [9:0] _T_2813 = {_T_2812[4'h0+:9], {{_T_2712}}};	// matmul/matmul-hw.mlir:12877:19, :12878:12, :12879:12, :12880:12
  wire [9:0] _T_2814 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12881:19, :12882:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12883:5
    if (rst)	// matmul/matmul-hw.mlir:12883:5
      _T_2811 <= _T_2814;	// matmul/matmul-hw.mlir:12886:7
    else	// matmul/matmul-hw.mlir:12883:5
      _T_2811 <= _T_2813;	// matmul/matmul-hw.mlir:12884:7
  end // always @(posedge)
  wire [9:0] _T_2816 = _T_2815;	// matmul/matmul-hw.mlir:12891:12
  wire [9:0] _T_2817 = {_T_2816[4'h0+:9], {{_T_2712}}};	// matmul/matmul-hw.mlir:12892:19, :12893:12, :12894:12, :12895:12
  wire [9:0] _T_2818 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12896:19, :12897:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12898:5
    if (rst)	// matmul/matmul-hw.mlir:12898:5
      _T_2815 <= _T_2818;	// matmul/matmul-hw.mlir:12901:7
    else	// matmul/matmul-hw.mlir:12898:5
      _T_2815 <= _T_2817;	// matmul/matmul-hw.mlir:12899:7
  end // always @(posedge)
  wire _T_2819 = _T_2815[4'h9];	// matmul/matmul-hw.mlir:12891:12, :12903:20, :12904:12
  assign _T_2142 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12905:12
  assign _T_2141 = _T_2819 ? A_p0_rd_data[4'h9] : 32'bx;	// matmul/matmul-hw.mlir:10176:19, :11112:15, :11113:12, :12906:12
  localparam [3:0] _T_2821 = 4'h0;	// matmul/matmul-hw.mlir:12909:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12910:5
    if (rst)	// matmul/matmul-hw.mlir:12910:5
      i_k_next_2820 <= _T_2821;	// matmul/matmul-hw.mlir:12913:7
    else	// matmul/matmul-hw.mlir:12910:5
      i_k_next_2820 <= i_k_next_2809;	// matmul/matmul-hw.mlir:12862:12, :12911:7
  end // always @(posedge)
  assign i_k_next_i_k_9 = i_k_next_2820;	// matmul/matmul-hw.mlir:12908:12, :12916:5
  //PROBE: i_k_next_i_k_9	// matmul/matmul-hw.mlir:12917:5
  assign _T_2140 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12918:12
  assign _T_2139 = _T_2819 ? i_k_next_2820 : 4'bx;	// matmul/matmul-hw.mlir:10174:18, :12908:12, :12919:12
  assign _T_2138 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12920:12
  wire [10:0] _T_2823 = _T_2822;	// matmul/matmul-hw.mlir:12922:12
  wire [10:0] _T_2824 = {_T_2823[4'h0+:10], {{_T_2712}}};	// matmul/matmul-hw.mlir:12923:19, :12924:12, :12925:12, :12926:12
  wire [10:0] _T_2825 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12927:19, :12928:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12929:5
    if (rst)	// matmul/matmul-hw.mlir:12929:5
      _T_2822 <= _T_2825;	// matmul/matmul-hw.mlir:12932:7
    else	// matmul/matmul-hw.mlir:12929:5
      _T_2822 <= _T_2824;	// matmul/matmul-hw.mlir:12930:7
  end // always @(posedge)
  wire [10:0] _T_2827 = _T_2826;	// matmul/matmul-hw.mlir:12937:12
  wire [10:0] _T_2828 = {_T_2827[4'h0+:10], {{_T_2712}}};	// matmul/matmul-hw.mlir:12938:19, :12939:12, :12940:12, :12941:12
  wire [10:0] _T_2829 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12942:19, :12943:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12944:5
    if (rst)	// matmul/matmul-hw.mlir:12944:5
      _T_2826 <= _T_2829;	// matmul/matmul-hw.mlir:12947:7
    else	// matmul/matmul-hw.mlir:12944:5
      _T_2826 <= _T_2828;	// matmul/matmul-hw.mlir:12945:7
  end // always @(posedge)
  wire _T_2830 = _T_2826[4'hA];	// matmul/matmul-hw.mlir:12937:12, :12949:20, :12950:12
  assign _T_2137 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12951:12
  assign _T_2136 = _T_2830 ? A_p0_rd_data[4'hA] : 32'bx;	// matmul/matmul-hw.mlir:10171:19, :11117:15, :11118:12, :12952:12
  localparam [3:0] _T_2832 = 4'h0;	// matmul/matmul-hw.mlir:12955:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12956:5
    if (rst)	// matmul/matmul-hw.mlir:12956:5
      i_k_next_2831 <= _T_2832;	// matmul/matmul-hw.mlir:12959:7
    else	// matmul/matmul-hw.mlir:12956:5
      i_k_next_2831 <= i_k_next_2820;	// matmul/matmul-hw.mlir:12908:12, :12957:7
  end // always @(posedge)
  assign i_k_next_i_k_10 = i_k_next_2831;	// matmul/matmul-hw.mlir:12954:12, :12962:5
  //PROBE: i_k_next_i_k_10	// matmul/matmul-hw.mlir:12963:5
  assign _T_2135 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12964:12
  assign _T_2134 = _T_2830 ? i_k_next_2831 : 4'bx;	// matmul/matmul-hw.mlir:10169:18, :12954:12, :12965:12
  assign _T_2133 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12966:12
  wire [11:0] _T_2834 = _T_2833;	// matmul/matmul-hw.mlir:12968:12
  wire [11:0] _T_2835 = {_T_2834[4'h0+:11], {{_T_2712}}};	// matmul/matmul-hw.mlir:12969:19, :12970:12, :12971:12, :12972:12
  wire [11:0] _T_2836 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12973:19, :12974:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12975:5
    if (rst)	// matmul/matmul-hw.mlir:12975:5
      _T_2833 <= _T_2836;	// matmul/matmul-hw.mlir:12978:7
    else	// matmul/matmul-hw.mlir:12975:5
      _T_2833 <= _T_2835;	// matmul/matmul-hw.mlir:12976:7
  end // always @(posedge)
  wire [11:0] _T_2838 = _T_2837;	// matmul/matmul-hw.mlir:12983:12
  wire [11:0] _T_2839 = {_T_2838[4'h0+:11], {{_T_2712}}};	// matmul/matmul-hw.mlir:12984:19, :12985:12, :12986:12, :12987:12
  wire [11:0] _T_2840 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:12988:19, :12989:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:12990:5
    if (rst)	// matmul/matmul-hw.mlir:12990:5
      _T_2837 <= _T_2840;	// matmul/matmul-hw.mlir:12993:7
    else	// matmul/matmul-hw.mlir:12990:5
      _T_2837 <= _T_2839;	// matmul/matmul-hw.mlir:12991:7
  end // always @(posedge)
  wire _T_2841 = _T_2837[4'hB];	// matmul/matmul-hw.mlir:12983:12, :12995:20, :12996:12
  assign _T_2132 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :12997:12
  assign _T_2131 = _T_2841 ? A_p0_rd_data[4'hB] : 32'bx;	// matmul/matmul-hw.mlir:10166:19, :11122:15, :11123:12, :12998:12
  localparam [3:0] _T_2843 = 4'h0;	// matmul/matmul-hw.mlir:13001:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13002:5
    if (rst)	// matmul/matmul-hw.mlir:13002:5
      i_k_next_2842 <= _T_2843;	// matmul/matmul-hw.mlir:13005:7
    else	// matmul/matmul-hw.mlir:13002:5
      i_k_next_2842 <= i_k_next_2831;	// matmul/matmul-hw.mlir:12954:12, :13003:7
  end // always @(posedge)
  assign i_k_next_i_k_11 = i_k_next_2842;	// matmul/matmul-hw.mlir:13000:12, :13008:5
  //PROBE: i_k_next_i_k_11	// matmul/matmul-hw.mlir:13009:5
  assign _T_2130 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13010:12
  assign _T_2129 = _T_2841 ? i_k_next_2842 : 4'bx;	// matmul/matmul-hw.mlir:10164:18, :13000:12, :13011:12
  assign _T_2128 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13012:12
  wire [12:0] _T_2845 = _T_2844;	// matmul/matmul-hw.mlir:13014:12
  wire [12:0] _T_2846 = {_T_2845[4'h0+:12], {{_T_2712}}};	// matmul/matmul-hw.mlir:13015:19, :13016:12, :13017:12, :13018:12
  wire [12:0] _T_2847 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13019:19, :13020:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13021:5
    if (rst)	// matmul/matmul-hw.mlir:13021:5
      _T_2844 <= _T_2847;	// matmul/matmul-hw.mlir:13024:7
    else	// matmul/matmul-hw.mlir:13021:5
      _T_2844 <= _T_2846;	// matmul/matmul-hw.mlir:13022:7
  end // always @(posedge)
  wire [12:0] _T_2849 = _T_2848;	// matmul/matmul-hw.mlir:13029:12
  wire [12:0] _T_2850 = {_T_2849[4'h0+:12], {{_T_2712}}};	// matmul/matmul-hw.mlir:13030:19, :13031:12, :13032:12, :13033:12
  wire [12:0] _T_2851 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13034:19, :13035:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13036:5
    if (rst)	// matmul/matmul-hw.mlir:13036:5
      _T_2848 <= _T_2851;	// matmul/matmul-hw.mlir:13039:7
    else	// matmul/matmul-hw.mlir:13036:5
      _T_2848 <= _T_2850;	// matmul/matmul-hw.mlir:13037:7
  end // always @(posedge)
  wire _T_2852 = _T_2848[4'hC];	// matmul/matmul-hw.mlir:13029:12, :13041:20, :13042:12
  assign _T_2127 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13043:12
  assign _T_2126 = _T_2852 ? A_p0_rd_data[4'hC] : 32'bx;	// matmul/matmul-hw.mlir:10161:19, :11127:15, :11128:12, :13044:12
  localparam [3:0] _T_2854 = 4'h0;	// matmul/matmul-hw.mlir:13047:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13048:5
    if (rst)	// matmul/matmul-hw.mlir:13048:5
      i_k_next_2853 <= _T_2854;	// matmul/matmul-hw.mlir:13051:7
    else	// matmul/matmul-hw.mlir:13048:5
      i_k_next_2853 <= i_k_next_2842;	// matmul/matmul-hw.mlir:13000:12, :13049:7
  end // always @(posedge)
  assign i_k_next_i_k_12 = i_k_next_2853;	// matmul/matmul-hw.mlir:13046:12, :13054:5
  //PROBE: i_k_next_i_k_12	// matmul/matmul-hw.mlir:13055:5
  assign _T_2125 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13056:12
  assign _T_2124 = _T_2852 ? i_k_next_2853 : 4'bx;	// matmul/matmul-hw.mlir:10159:18, :13046:12, :13057:12
  assign _T_2123 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13058:12
  wire [13:0] _T_2856 = _T_2855;	// matmul/matmul-hw.mlir:13060:12
  wire [13:0] _T_2857 = {_T_2856[4'h0+:13], {{_T_2712}}};	// matmul/matmul-hw.mlir:13061:19, :13062:12, :13063:12, :13064:12
  wire [13:0] _T_2858 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13065:19, :13066:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13067:5
    if (rst)	// matmul/matmul-hw.mlir:13067:5
      _T_2855 <= _T_2858;	// matmul/matmul-hw.mlir:13070:7
    else	// matmul/matmul-hw.mlir:13067:5
      _T_2855 <= _T_2857;	// matmul/matmul-hw.mlir:13068:7
  end // always @(posedge)
  wire [13:0] _T_2860 = _T_2859;	// matmul/matmul-hw.mlir:13075:12
  wire [13:0] _T_2861 = {_T_2860[4'h0+:13], {{_T_2712}}};	// matmul/matmul-hw.mlir:13076:19, :13077:12, :13078:12, :13079:12
  wire [13:0] _T_2862 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13080:19, :13081:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13082:5
    if (rst)	// matmul/matmul-hw.mlir:13082:5
      _T_2859 <= _T_2862;	// matmul/matmul-hw.mlir:13085:7
    else	// matmul/matmul-hw.mlir:13082:5
      _T_2859 <= _T_2861;	// matmul/matmul-hw.mlir:13083:7
  end // always @(posedge)
  wire _T_2863 = _T_2859[4'hD];	// matmul/matmul-hw.mlir:13075:12, :13087:20, :13088:12
  assign _T_2122 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13089:12
  assign _T_2121 = _T_2863 ? A_p0_rd_data[4'hD] : 32'bx;	// matmul/matmul-hw.mlir:10156:19, :11132:15, :11133:12, :13090:12
  localparam [3:0] _T_2865 = 4'h0;	// matmul/matmul-hw.mlir:13093:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13094:5
    if (rst)	// matmul/matmul-hw.mlir:13094:5
      i_k_next_2864 <= _T_2865;	// matmul/matmul-hw.mlir:13097:7
    else	// matmul/matmul-hw.mlir:13094:5
      i_k_next_2864 <= i_k_next_2853;	// matmul/matmul-hw.mlir:13046:12, :13095:7
  end // always @(posedge)
  assign i_k_next_i_k_13 = i_k_next_2864;	// matmul/matmul-hw.mlir:13092:12, :13100:5
  //PROBE: i_k_next_i_k_13	// matmul/matmul-hw.mlir:13101:5
  assign _T_2120 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13102:12
  assign _T_2119 = _T_2863 ? i_k_next_2864 : 4'bx;	// matmul/matmul-hw.mlir:10154:18, :13092:12, :13103:12
  assign _T_2118 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13104:12
  wire [14:0] _T_2867 = _T_2866;	// matmul/matmul-hw.mlir:13106:12
  wire [14:0] _T_2868 = {_T_2867[4'h0+:14], {{_T_2712}}};	// matmul/matmul-hw.mlir:13107:19, :13108:12, :13109:12, :13110:12
  wire [14:0] _T_2869 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13111:19, :13112:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13113:5
    if (rst)	// matmul/matmul-hw.mlir:13113:5
      _T_2866 <= _T_2869;	// matmul/matmul-hw.mlir:13116:7
    else	// matmul/matmul-hw.mlir:13113:5
      _T_2866 <= _T_2868;	// matmul/matmul-hw.mlir:13114:7
  end // always @(posedge)
  wire [14:0] _T_2871 = _T_2870;	// matmul/matmul-hw.mlir:13121:12
  wire [14:0] _T_2872 = {_T_2871[4'h0+:14], {{_T_2712}}};	// matmul/matmul-hw.mlir:13122:19, :13123:12, :13124:12, :13125:12
  wire [14:0] _T_2873 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13126:19, :13127:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13128:5
    if (rst)	// matmul/matmul-hw.mlir:13128:5
      _T_2870 <= _T_2873;	// matmul/matmul-hw.mlir:13131:7
    else	// matmul/matmul-hw.mlir:13128:5
      _T_2870 <= _T_2872;	// matmul/matmul-hw.mlir:13129:7
  end // always @(posedge)
  wire _T_2874 = _T_2870[4'hE];	// matmul/matmul-hw.mlir:13121:12, :13133:20, :13134:12
  assign _T_2117 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13135:12
  assign _T_2116 = _T_2874 ? A_p0_rd_data[4'hE] : 32'bx;	// matmul/matmul-hw.mlir:10151:19, :11137:15, :11138:12, :13136:12
  localparam [3:0] _T_2876 = 4'h0;	// matmul/matmul-hw.mlir:13139:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13140:5
    if (rst)	// matmul/matmul-hw.mlir:13140:5
      i_k_next_2875 <= _T_2876;	// matmul/matmul-hw.mlir:13143:7
    else	// matmul/matmul-hw.mlir:13140:5
      i_k_next_2875 <= i_k_next_2864;	// matmul/matmul-hw.mlir:13092:12, :13141:7
  end // always @(posedge)
  assign i_k_next_i_k_14 = i_k_next_2875;	// matmul/matmul-hw.mlir:13138:12, :13146:5
  //PROBE: i_k_next_i_k_14	// matmul/matmul-hw.mlir:13147:5
  assign _T_2115 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13148:12
  assign _T_2114 = _T_2874 ? i_k_next_2875 : 4'bx;	// matmul/matmul-hw.mlir:10149:18, :13138:12, :13149:12
  assign _T_2113 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13150:12
  wire [15:0] _T_2878 = _T_2877;	// matmul/matmul-hw.mlir:13152:12
  wire [15:0] _T_2879 = {_T_2878[4'h0+:15], {{_T_2712}}};	// matmul/matmul-hw.mlir:13153:19, :13154:12, :13155:12, :13156:12
  wire [15:0] _T_2880 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13157:19, :13158:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13159:5
    if (rst)	// matmul/matmul-hw.mlir:13159:5
      _T_2877 <= _T_2880;	// matmul/matmul-hw.mlir:13162:7
    else	// matmul/matmul-hw.mlir:13159:5
      _T_2877 <= _T_2879;	// matmul/matmul-hw.mlir:13160:7
  end // always @(posedge)
  wire [15:0] _T_2882 = _T_2881;	// matmul/matmul-hw.mlir:13167:12
  wire [15:0] _T_2883 = {_T_2882[4'h0+:15], {{_T_2712}}};	// matmul/matmul-hw.mlir:13168:19, :13169:12, :13170:12, :13171:12
  wire [15:0] _T_2884 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13172:19, :13173:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13174:5
    if (rst)	// matmul/matmul-hw.mlir:13174:5
      _T_2881 <= _T_2884;	// matmul/matmul-hw.mlir:13177:7
    else	// matmul/matmul-hw.mlir:13174:5
      _T_2881 <= _T_2883;	// matmul/matmul-hw.mlir:13175:7
  end // always @(posedge)
  wire _T_2885 = _T_2881[4'hF];	// matmul/matmul-hw.mlir:13167:12, :13179:20, :13180:12
  assign _T_2112 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13181:12
  assign _T_2111 = _T_2885 ? A_p0_rd_data[4'hF] : 32'bx;	// matmul/matmul-hw.mlir:10146:19, :11142:15, :11143:12, :13182:12
  localparam [3:0] _T_2887 = 4'h0;	// matmul/matmul-hw.mlir:13185:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13186:5
    if (rst)	// matmul/matmul-hw.mlir:13186:5
      i_k_next_2886 <= _T_2887;	// matmul/matmul-hw.mlir:13189:7
    else	// matmul/matmul-hw.mlir:13186:5
      i_k_next_2886 <= i_k_next_2875;	// matmul/matmul-hw.mlir:13138:12, :13187:7
  end // always @(posedge)
  assign i_k_next_i_k_15 = i_k_next_2886;	// matmul/matmul-hw.mlir:13184:12, :13192:5
  //PROBE: i_k_next_i_k_15	// matmul/matmul-hw.mlir:13193:5
  assign _T_2110 = _T_2731 ? 1'h1 : _T_1388;	// matmul/matmul-hw.mlir:8029:13, :13194:12, :14226:13
  assign _T_2109 = _T_2731 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13195:12
  assign _T_2108 = _T_2731 ? A_reg_bank0_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10143:19, :12215:31, :13196:12
  assign _T_2107 = _T_2742 ? 1'h1 : _T_1383;	// matmul/matmul-hw.mlir:8029:13, :13197:12, :14248:13
  assign _T_2106 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13198:12
  assign _T_2105 = _T_2742 ? A_reg_bank1_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10140:19, :12216:31, :13199:12
  assign _T_2104 = _T_2753 ? 1'h1 : _T_1378;	// matmul/matmul-hw.mlir:8029:13, :13200:12, :14270:13
  assign _T_2103 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13201:12
  assign _T_2102 = _T_2753 ? A_reg_bank2_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10137:19, :12217:31, :13202:12
  assign _T_2101 = _T_2764 ? 1'h1 : _T_1373;	// matmul/matmul-hw.mlir:8029:13, :13203:12, :14292:13
  assign _T_2100 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13204:12
  assign _T_2099 = _T_2764 ? A_reg_bank3_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10134:19, :12218:31, :13205:12
  assign _T_2098 = _T_2775 ? 1'h1 : _T_1368;	// matmul/matmul-hw.mlir:8029:13, :13206:12, :14314:13
  assign _T_2097 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13207:12
  assign _T_2096 = _T_2775 ? A_reg_bank4_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10131:19, :12219:31, :13208:12
  assign _T_2095 = _T_2786 ? 1'h1 : _T_1363;	// matmul/matmul-hw.mlir:8029:13, :13209:12, :14336:13
  assign _T_2094 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13210:12
  assign _T_2093 = _T_2786 ? A_reg_bank5_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10128:19, :12220:31, :13211:12
  assign _T_2092 = _T_2797 ? 1'h1 : _T_1358;	// matmul/matmul-hw.mlir:8029:13, :13212:12, :14358:13
  assign _T_2091 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13213:12
  assign _T_2090 = _T_2797 ? A_reg_bank6_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10125:19, :12221:31, :13214:12
  assign _T_2089 = _T_2808 ? 1'h1 : _T_1353;	// matmul/matmul-hw.mlir:8029:13, :13215:12, :14380:13
  assign _T_2088 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13216:12
  assign _T_2087 = _T_2808 ? A_reg_bank7_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10122:19, :12222:31, :13217:12
  assign _T_2086 = _T_2819 ? 1'h1 : _T_1348;	// matmul/matmul-hw.mlir:8029:13, :13218:12, :14402:13
  assign _T_2085 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13219:12
  assign _T_2084 = _T_2819 ? A_reg_bank8_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10119:19, :12223:31, :13220:12
  assign _T_2083 = _T_2830 ? 1'h1 : _T_1343;	// matmul/matmul-hw.mlir:8029:13, :13221:12, :14424:13
  assign _T_2082 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13222:12
  assign _T_2081 = _T_2830 ? A_reg_bank9_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10116:19, :12224:31, :13223:12
  assign _T_2080 = _T_2841 ? 1'h1 : _T_1338;	// matmul/matmul-hw.mlir:8029:13, :13224:12, :14446:13
  assign _T_2079 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13225:12
  assign _T_2078 = _T_2841 ? A_reg_bank10_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10113:19, :12225:32, :13226:12
  assign _T_2077 = _T_2852 ? 1'h1 : _T_1333;	// matmul/matmul-hw.mlir:8029:13, :13227:12, :14468:13
  assign _T_2076 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13228:12
  assign _T_2075 = _T_2852 ? A_reg_bank11_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10110:19, :12226:32, :13229:12
  assign _T_2074 = _T_2863 ? 1'h1 : _T_1328;	// matmul/matmul-hw.mlir:8029:13, :13230:12, :14490:13
  assign _T_2073 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13231:12
  assign _T_2072 = _T_2863 ? A_reg_bank12_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10107:19, :12227:32, :13232:12
  assign _T_2071 = _T_2874 ? 1'h1 : _T_1323;	// matmul/matmul-hw.mlir:8029:13, :13233:12, :14512:13
  assign _T_2070 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13234:12
  assign _T_2069 = _T_2874 ? A_reg_bank13_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10104:19, :12228:32, :13235:12
  assign _T_2068 = _T_2885 ? 1'h1 : _T_1318;	// matmul/matmul-hw.mlir:8029:13, :13236:12, :14534:13
  assign _T_2067 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13237:12
  assign _T_2066 = _T_2885 ? A_reg_bank14_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10101:19, :12229:32, :13238:12
  wire [16:0] _T_2889 = _T_2888;	// matmul/matmul-hw.mlir:13240:12
  wire [16:0] _T_2890 = {_T_2889[5'h0+:16], {{_T_2712}}};	// matmul/matmul-hw.mlir:13241:14, :13242:12, :13243:12, :13244:12
  wire [16:0] _T_2891 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13245:19, :13246:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13247:5
    if (rst)	// matmul/matmul-hw.mlir:13247:5
      _T_2888 <= _T_2891;	// matmul/matmul-hw.mlir:13250:7
    else	// matmul/matmul-hw.mlir:13247:5
      _T_2888 <= _T_2890;	// matmul/matmul-hw.mlir:13248:7
  end // always @(posedge)
  wire _T_2892 = _T_2888[5'h10];	// matmul/matmul-hw.mlir:13240:12, :13252:16, :13253:12
  assign _T_2065 = _T_2892 ? 1'h1 : _T_1313;	// matmul/matmul-hw.mlir:8029:13, :13254:12, :14556:13
  assign _T_2064 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13255:12
  assign _T_2063 = _T_2892 ? A_reg_bank15_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10098:19, :12230:32, :13256:12
  assign _T_2062 = _T_2742 ? 1'h1 : _T_1301;	// matmul/matmul-hw.mlir:8029:13, :13257:12, :14693:13
  assign _T_2061 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13258:12
  assign _T_2060 = _T_2742 ? A_reg_bank16_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10095:19, :12231:32, :13259:12
  assign _T_2059 = _T_2753 ? 1'h1 : _T_1296;	// matmul/matmul-hw.mlir:8029:13, :13260:12, :14723:13
  assign _T_2058 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13261:12
  assign _T_2057 = _T_2753 ? A_reg_bank17_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10092:19, :12232:32, :13262:12
  assign _T_2056 = _T_2764 ? 1'h1 : _T_1291;	// matmul/matmul-hw.mlir:8029:13, :13263:12, :14753:13
  assign _T_2055 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13264:12
  assign _T_2054 = _T_2764 ? A_reg_bank18_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10089:19, :12233:32, :13265:12
  assign _T_2053 = _T_2775 ? 1'h1 : _T_1286;	// matmul/matmul-hw.mlir:8029:13, :13266:12, :14783:13
  assign _T_2052 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13267:12
  assign _T_2051 = _T_2775 ? A_reg_bank19_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10086:19, :12234:32, :13268:12
  assign _T_2050 = _T_2786 ? 1'h1 : _T_1281;	// matmul/matmul-hw.mlir:8029:13, :13269:12, :14813:13
  assign _T_2049 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13270:12
  assign _T_2048 = _T_2786 ? A_reg_bank20_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10083:19, :12235:32, :13271:12
  assign _T_2047 = _T_2797 ? 1'h1 : _T_1276;	// matmul/matmul-hw.mlir:8029:13, :13272:12, :14843:13
  assign _T_2046 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13273:12
  assign _T_2045 = _T_2797 ? A_reg_bank21_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10080:19, :12236:32, :13274:12
  assign _T_2044 = _T_2808 ? 1'h1 : _T_1271;	// matmul/matmul-hw.mlir:8029:13, :13275:12, :14873:13
  assign _T_2043 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13276:12
  assign _T_2042 = _T_2808 ? A_reg_bank22_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10077:19, :12237:32, :13277:12
  assign _T_2041 = _T_2819 ? 1'h1 : _T_1266;	// matmul/matmul-hw.mlir:8029:13, :13278:12, :14903:13
  assign _T_2040 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13279:12
  assign _T_2039 = _T_2819 ? A_reg_bank23_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10074:19, :12238:32, :13280:12
  assign _T_2038 = _T_2830 ? 1'h1 : _T_1261;	// matmul/matmul-hw.mlir:8029:13, :13281:12, :14933:13
  assign _T_2037 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13282:12
  assign _T_2036 = _T_2830 ? A_reg_bank24_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10071:19, :12239:32, :13283:12
  assign _T_2035 = _T_2841 ? 1'h1 : _T_1256;	// matmul/matmul-hw.mlir:8029:13, :13284:12, :14963:13
  assign _T_2034 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13285:12
  assign _T_2033 = _T_2841 ? A_reg_bank25_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10068:19, :12240:32, :13286:12
  assign _T_2032 = _T_2852 ? 1'h1 : _T_1251;	// matmul/matmul-hw.mlir:8029:13, :13287:12, :14993:13
  assign _T_2031 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13288:12
  assign _T_2030 = _T_2852 ? A_reg_bank26_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10065:19, :12241:32, :13289:12
  assign _T_2029 = _T_2863 ? 1'h1 : _T_1246;	// matmul/matmul-hw.mlir:8029:13, :13290:12, :15023:13
  assign _T_2028 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13291:12
  assign _T_2027 = _T_2863 ? A_reg_bank27_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10062:19, :12242:32, :13292:12
  assign _T_2026 = _T_2874 ? 1'h1 : _T_1241;	// matmul/matmul-hw.mlir:8029:13, :13293:12, :15053:13
  assign _T_2025 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13294:12
  assign _T_2024 = _T_2874 ? A_reg_bank28_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10059:19, :12243:32, :13295:12
  assign _T_2023 = _T_2885 ? 1'h1 : _T_1236;	// matmul/matmul-hw.mlir:8029:13, :13296:12, :15083:13
  assign _T_2022 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13297:12
  assign _T_2021 = _T_2885 ? A_reg_bank29_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10056:19, :12244:32, :13298:12
  assign _T_2020 = _T_2892 ? 1'h1 : _T_1231;	// matmul/matmul-hw.mlir:8029:13, :13299:12, :15113:13
  assign _T_2019 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13300:12
  assign _T_2018 = _T_2892 ? A_reg_bank30_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10053:19, :12245:32, :13301:12
  wire [17:0] _T_2894 = _T_2893;	// matmul/matmul-hw.mlir:13303:12
  wire [17:0] _T_2895 = {_T_2894[5'h0+:17], {{_T_2712}}};	// matmul/matmul-hw.mlir:13304:19, :13305:12, :13306:12, :13307:12
  wire [17:0] _T_2896 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13308:19, :13309:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13310:5
    if (rst)	// matmul/matmul-hw.mlir:13310:5
      _T_2893 <= _T_2896;	// matmul/matmul-hw.mlir:13313:7
    else	// matmul/matmul-hw.mlir:13310:5
      _T_2893 <= _T_2895;	// matmul/matmul-hw.mlir:13311:7
  end // always @(posedge)
  wire _T_2897 = _T_2893[5'h11];	// matmul/matmul-hw.mlir:13303:12, :13315:16, :13316:12
  assign _T_2017 = _T_2897 ? 1'h1 : _T_1226;	// matmul/matmul-hw.mlir:8029:13, :13317:12, :15143:13
  assign _T_2016 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13318:12
  assign _T_2015 = _T_2897 ? A_reg_bank31_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10050:19, :12246:32, :13319:12
  assign _T_2014 = _T_2753 ? 1'h1 : _T_1214;	// matmul/matmul-hw.mlir:8029:13, :13320:12, :15288:13
  assign _T_2013 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13321:12
  assign _T_2012 = _T_2753 ? A_reg_bank32_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10047:19, :12247:32, :13322:12
  assign _T_2011 = _T_2764 ? 1'h1 : _T_1209;	// matmul/matmul-hw.mlir:8029:13, :13323:12, :15318:13
  assign _T_2010 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13324:12
  assign _T_2009 = _T_2764 ? A_reg_bank33_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10044:19, :12248:32, :13325:12
  assign _T_2008 = _T_2775 ? 1'h1 : _T_1204;	// matmul/matmul-hw.mlir:8029:13, :13326:12, :15348:13
  assign _T_2007 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13327:12
  assign _T_2006 = _T_2775 ? A_reg_bank34_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10041:19, :12249:32, :13328:12
  assign _T_2005 = _T_2786 ? 1'h1 : _T_1199;	// matmul/matmul-hw.mlir:8029:13, :13329:12, :15378:13
  assign _T_2004 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13330:12
  assign _T_2003 = _T_2786 ? A_reg_bank35_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10038:19, :12250:32, :13331:12
  assign _T_2002 = _T_2797 ? 1'h1 : _T_1194;	// matmul/matmul-hw.mlir:8029:13, :13332:12, :15408:13
  assign _T_2001 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13333:12
  assign _T_2000 = _T_2797 ? A_reg_bank36_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10035:19, :12251:32, :13334:12
  assign _T_1999 = _T_2808 ? 1'h1 : _T_1189;	// matmul/matmul-hw.mlir:8029:13, :13335:12, :15438:13
  assign _T_1998 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13336:12
  assign _T_1997 = _T_2808 ? A_reg_bank37_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10032:19, :12252:32, :13337:12
  assign _T_1996 = _T_2819 ? 1'h1 : _T_1184;	// matmul/matmul-hw.mlir:8029:13, :13338:12, :15468:13
  assign _T_1995 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13339:12
  assign _T_1994 = _T_2819 ? A_reg_bank38_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10029:19, :12253:32, :13340:12
  assign _T_1993 = _T_2830 ? 1'h1 : _T_1179;	// matmul/matmul-hw.mlir:8029:13, :13341:12, :15498:13
  assign _T_1992 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13342:12
  assign _T_1991 = _T_2830 ? A_reg_bank39_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10026:19, :12254:32, :13343:12
  assign _T_1990 = _T_2841 ? 1'h1 : _T_1174;	// matmul/matmul-hw.mlir:8029:13, :13344:12, :15528:13
  assign _T_1989 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13345:12
  assign _T_1988 = _T_2841 ? A_reg_bank40_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10023:19, :12255:32, :13346:12
  assign _T_1987 = _T_2852 ? 1'h1 : _T_1169;	// matmul/matmul-hw.mlir:8029:13, :13347:12, :15558:13
  assign _T_1986 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13348:12
  assign _T_1985 = _T_2852 ? A_reg_bank41_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10020:19, :12256:32, :13349:12
  assign _T_1984 = _T_2863 ? 1'h1 : _T_1164;	// matmul/matmul-hw.mlir:8029:13, :13350:12, :15588:13
  assign _T_1983 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13351:12
  assign _T_1982 = _T_2863 ? A_reg_bank42_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10017:19, :12257:32, :13352:12
  assign _T_1981 = _T_2874 ? 1'h1 : _T_1159;	// matmul/matmul-hw.mlir:8029:13, :13353:12, :15618:13
  assign _T_1980 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13354:12
  assign _T_1979 = _T_2874 ? A_reg_bank43_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10014:19, :12258:32, :13355:12
  assign _T_1978 = _T_2885 ? 1'h1 : _T_1154;	// matmul/matmul-hw.mlir:8029:13, :13356:12, :15648:13
  assign _T_1977 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13357:12
  assign _T_1976 = _T_2885 ? A_reg_bank44_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10011:19, :12259:32, :13358:12
  assign _T_1975 = _T_2892 ? 1'h1 : _T_1149;	// matmul/matmul-hw.mlir:8029:13, :13359:12, :15678:13
  assign _T_1974 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13360:12
  assign _T_1973 = _T_2892 ? A_reg_bank45_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10008:19, :12260:32, :13361:12
  assign _T_1972 = _T_2897 ? 1'h1 : _T_1144;	// matmul/matmul-hw.mlir:8029:13, :13362:12, :15708:13
  assign _T_1971 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13363:12
  assign _T_1970 = _T_2897 ? A_reg_bank46_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10005:19, :12261:32, :13364:12
  wire [18:0] _T_2899 = _T_2898;	// matmul/matmul-hw.mlir:13366:12
  wire [18:0] _T_2900 = {_T_2899[5'h0+:18], {{_T_2712}}};	// matmul/matmul-hw.mlir:13367:19, :13368:12, :13369:12, :13370:12
  wire [18:0] _T_2901 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13371:19, :13372:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13373:5
    if (rst)	// matmul/matmul-hw.mlir:13373:5
      _T_2898 <= _T_2901;	// matmul/matmul-hw.mlir:13376:7
    else	// matmul/matmul-hw.mlir:13373:5
      _T_2898 <= _T_2900;	// matmul/matmul-hw.mlir:13374:7
  end // always @(posedge)
  wire _T_2902 = _T_2898[5'h12];	// matmul/matmul-hw.mlir:13366:12, :13378:16, :13379:12
  assign _T_1969 = _T_2902 ? 1'h1 : _T_1139;	// matmul/matmul-hw.mlir:8029:13, :13380:12, :15738:13
  assign _T_1968 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13381:12
  assign _T_1967 = _T_2902 ? A_reg_bank47_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:10002:19, :12262:32, :13382:12
  assign _T_1966 = _T_2764 ? 1'h1 : _T_1127;	// matmul/matmul-hw.mlir:8029:13, :13383:12, :15883:13
  assign _T_1965 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13384:12
  assign _T_1964 = _T_2764 ? A_reg_bank48_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9999:19, :12263:32, :13385:12
  assign _T_1963 = _T_2775 ? 1'h1 : _T_1122;	// matmul/matmul-hw.mlir:8029:13, :13386:12, :15913:13
  assign _T_1962 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13387:12
  assign _T_1961 = _T_2775 ? A_reg_bank49_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9996:19, :12264:32, :13388:12
  assign _T_1960 = _T_2786 ? 1'h1 : _T_1117;	// matmul/matmul-hw.mlir:8029:13, :13389:12, :15943:13
  assign _T_1959 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13390:12
  assign _T_1958 = _T_2786 ? A_reg_bank50_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9993:19, :12265:32, :13391:12
  assign _T_1957 = _T_2797 ? 1'h1 : _T_1112;	// matmul/matmul-hw.mlir:8029:13, :13392:12, :15973:13
  assign _T_1956 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13393:12
  assign _T_1955 = _T_2797 ? A_reg_bank51_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9990:19, :12266:32, :13394:12
  assign _T_1954 = _T_2808 ? 1'h1 : _T_1107;	// matmul/matmul-hw.mlir:8029:13, :13395:12, :16003:13
  assign _T_1953 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13396:12
  assign _T_1952 = _T_2808 ? A_reg_bank52_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9987:19, :12267:32, :13397:12
  assign _T_1951 = _T_2819 ? 1'h1 : _T_1102;	// matmul/matmul-hw.mlir:8029:13, :13398:12, :16033:13
  assign _T_1950 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13399:12
  assign _T_1949 = _T_2819 ? A_reg_bank53_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9984:19, :12268:32, :13400:12
  assign _T_1948 = _T_2830 ? 1'h1 : _T_1097;	// matmul/matmul-hw.mlir:8029:13, :13401:12, :16063:13
  assign _T_1947 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13402:12
  assign _T_1946 = _T_2830 ? A_reg_bank54_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9981:19, :12269:32, :13403:12
  assign _T_1945 = _T_2841 ? 1'h1 : _T_1092;	// matmul/matmul-hw.mlir:8029:13, :13404:12, :16093:13
  assign _T_1944 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13405:12
  assign _T_1943 = _T_2841 ? A_reg_bank55_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9978:19, :12270:32, :13406:12
  assign _T_1942 = _T_2852 ? 1'h1 : _T_1087;	// matmul/matmul-hw.mlir:8029:13, :13407:12, :16123:13
  assign _T_1941 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13408:12
  assign _T_1940 = _T_2852 ? A_reg_bank56_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9975:19, :12271:32, :13409:12
  assign _T_1939 = _T_2863 ? 1'h1 : _T_1082;	// matmul/matmul-hw.mlir:8029:13, :13410:12, :16153:13
  assign _T_1938 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13411:12
  assign _T_1937 = _T_2863 ? A_reg_bank57_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9972:19, :12272:32, :13412:12
  assign _T_1936 = _T_2874 ? 1'h1 : _T_1077;	// matmul/matmul-hw.mlir:8029:13, :13413:12, :16183:13
  assign _T_1935 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13414:12
  assign _T_1934 = _T_2874 ? A_reg_bank58_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9969:19, :12273:32, :13415:12
  assign _T_1933 = _T_2885 ? 1'h1 : _T_1072;	// matmul/matmul-hw.mlir:8029:13, :13416:12, :16213:13
  assign _T_1932 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13417:12
  assign _T_1931 = _T_2885 ? A_reg_bank59_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9966:19, :12274:32, :13418:12
  assign _T_1930 = _T_2892 ? 1'h1 : _T_1067;	// matmul/matmul-hw.mlir:8029:13, :13419:12, :16243:13
  assign _T_1929 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13420:12
  assign _T_1928 = _T_2892 ? A_reg_bank60_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9963:19, :12275:32, :13421:12
  assign _T_1927 = _T_2897 ? 1'h1 : _T_1062;	// matmul/matmul-hw.mlir:8029:13, :13422:12, :16273:13
  assign _T_1926 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13423:12
  assign _T_1925 = _T_2897 ? A_reg_bank61_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9960:19, :12276:32, :13424:12
  assign _T_1924 = _T_2902 ? 1'h1 : _T_1057;	// matmul/matmul-hw.mlir:8029:13, :13425:12, :16303:13
  assign _T_1923 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13426:12
  assign _T_1922 = _T_2902 ? A_reg_bank62_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9957:19, :12277:32, :13427:12
  wire [19:0] _T_2904 = _T_2903;	// matmul/matmul-hw.mlir:13429:12
  wire [19:0] _T_2905 = {_T_2904[5'h0+:19], {{_T_2712}}};	// matmul/matmul-hw.mlir:13430:19, :13431:12, :13432:12, :13433:12
  wire [19:0] _T_2906 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13434:19, :13435:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13436:5
    if (rst)	// matmul/matmul-hw.mlir:13436:5
      _T_2903 <= _T_2906;	// matmul/matmul-hw.mlir:13439:7
    else	// matmul/matmul-hw.mlir:13436:5
      _T_2903 <= _T_2905;	// matmul/matmul-hw.mlir:13437:7
  end // always @(posedge)
  wire _T_2907 = _T_2903[5'h13];	// matmul/matmul-hw.mlir:13429:12, :13441:16, :13442:12
  assign _T_1921 = _T_2907 ? 1'h1 : _T_1052;	// matmul/matmul-hw.mlir:8029:13, :13443:12, :16333:13
  assign _T_1920 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13444:12
  assign _T_1919 = _T_2907 ? A_reg_bank63_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9954:19, :12278:32, :13445:12
  assign _T_1918 = _T_2775 ? 1'h1 : _T_1040;	// matmul/matmul-hw.mlir:8029:13, :13446:12, :16478:13
  assign _T_1917 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13447:12
  assign _T_1916 = _T_2775 ? A_reg_bank64_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9951:19, :12279:32, :13448:12
  assign _T_1915 = _T_2786 ? 1'h1 : _T_1035;	// matmul/matmul-hw.mlir:8029:13, :13449:12, :16508:13
  assign _T_1914 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13450:12
  assign _T_1913 = _T_2786 ? A_reg_bank65_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9948:19, :12280:32, :13451:12
  assign _T_1912 = _T_2797 ? 1'h1 : _T_1030;	// matmul/matmul-hw.mlir:8029:13, :13452:12, :16538:13
  assign _T_1911 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13453:12
  assign _T_1910 = _T_2797 ? A_reg_bank66_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9945:19, :12281:32, :13454:12
  assign _T_1909 = _T_2808 ? 1'h1 : _T_1025;	// matmul/matmul-hw.mlir:8029:13, :13455:12, :16568:13
  assign _T_1908 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13456:12
  assign _T_1907 = _T_2808 ? A_reg_bank67_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9942:19, :12282:32, :13457:12
  assign _T_1906 = _T_2819 ? 1'h1 : _T_1020;	// matmul/matmul-hw.mlir:8029:13, :13458:12, :16598:13
  assign _T_1905 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13459:12
  assign _T_1904 = _T_2819 ? A_reg_bank68_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9939:19, :12283:32, :13460:12
  assign _T_1903 = _T_2830 ? 1'h1 : _T_1015;	// matmul/matmul-hw.mlir:8029:13, :13461:12, :16628:13
  assign _T_1902 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13462:12
  assign _T_1901 = _T_2830 ? A_reg_bank69_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9936:19, :12284:32, :13463:12
  assign _T_1900 = _T_2841 ? 1'h1 : _T_1010;	// matmul/matmul-hw.mlir:8029:13, :13464:12, :16658:13
  assign _T_1899 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13465:12
  assign _T_1898 = _T_2841 ? A_reg_bank70_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9933:19, :12285:32, :13466:12
  assign _T_1897 = _T_2852 ? 1'h1 : _T_1005;	// matmul/matmul-hw.mlir:8029:13, :13467:12, :16688:13
  assign _T_1896 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13468:12
  assign _T_1895 = _T_2852 ? A_reg_bank71_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9930:19, :12286:32, :13469:12
  assign _T_1894 = _T_2863 ? 1'h1 : _T_1000;	// matmul/matmul-hw.mlir:8029:13, :13470:12, :16718:13
  assign _T_1893 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13471:12
  assign _T_1892 = _T_2863 ? A_reg_bank72_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9927:19, :12287:32, :13472:12
  assign _T_1891 = _T_2874 ? 1'h1 : _T_995;	// matmul/matmul-hw.mlir:8029:13, :13473:12, :16748:13
  assign _T_1890 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13474:12
  assign _T_1889 = _T_2874 ? A_reg_bank73_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9924:19, :12288:32, :13475:12
  assign _T_1888 = _T_2885 ? 1'h1 : _T_990;	// matmul/matmul-hw.mlir:8029:13, :13476:12, :16778:13
  assign _T_1887 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13477:12
  assign _T_1886 = _T_2885 ? A_reg_bank74_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9921:19, :12289:32, :13478:12
  assign _T_1885 = _T_2892 ? 1'h1 : _T_985;	// matmul/matmul-hw.mlir:8029:13, :13479:12, :16808:13
  assign _T_1884 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13480:12
  assign _T_1883 = _T_2892 ? A_reg_bank75_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9918:19, :12290:32, :13481:12
  assign _T_1882 = _T_2897 ? 1'h1 : _T_980;	// matmul/matmul-hw.mlir:8029:13, :13482:12, :16838:13
  assign _T_1881 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13483:12
  assign _T_1880 = _T_2897 ? A_reg_bank76_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9915:19, :12291:32, :13484:12
  assign _T_1879 = _T_2902 ? 1'h1 : _T_975;	// matmul/matmul-hw.mlir:8029:13, :13485:12, :16868:13
  assign _T_1878 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13486:12
  assign _T_1877 = _T_2902 ? A_reg_bank77_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9912:19, :12292:32, :13487:12
  assign _T_1876 = _T_2907 ? 1'h1 : _T_970;	// matmul/matmul-hw.mlir:8029:13, :13488:12, :16898:13
  assign _T_1875 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13489:12
  assign _T_1874 = _T_2907 ? A_reg_bank78_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9909:19, :12293:32, :13490:12
  wire [20:0] _T_2909 = _T_2908;	// matmul/matmul-hw.mlir:13492:12
  wire [20:0] _T_2910 = {_T_2909[5'h0+:20], {{_T_2712}}};	// matmul/matmul-hw.mlir:13493:19, :13494:12, :13495:12, :13496:12
  wire [20:0] _T_2911 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13497:19, :13498:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13499:5
    if (rst)	// matmul/matmul-hw.mlir:13499:5
      _T_2908 <= _T_2911;	// matmul/matmul-hw.mlir:13502:7
    else	// matmul/matmul-hw.mlir:13499:5
      _T_2908 <= _T_2910;	// matmul/matmul-hw.mlir:13500:7
  end // always @(posedge)
  wire _T_2912 = _T_2908[5'h14];	// matmul/matmul-hw.mlir:13492:12, :13504:16, :13505:12
  assign _T_1873 = _T_2912 ? 1'h1 : _T_965;	// matmul/matmul-hw.mlir:8029:13, :13506:12, :16928:13
  assign _T_1872 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13507:12
  assign _T_1871 = _T_2912 ? A_reg_bank79_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9906:19, :12294:32, :13508:12
  assign _T_1870 = _T_2786 ? 1'h1 : _T_953;	// matmul/matmul-hw.mlir:8029:13, :13509:12, :17073:13
  assign _T_1869 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13510:12
  assign _T_1868 = _T_2786 ? A_reg_bank80_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9903:19, :12295:32, :13511:12
  assign _T_1867 = _T_2797 ? 1'h1 : _T_948;	// matmul/matmul-hw.mlir:8029:13, :13512:12, :17103:13
  assign _T_1866 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13513:12
  assign _T_1865 = _T_2797 ? A_reg_bank81_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9900:19, :12296:32, :13514:12
  assign _T_1864 = _T_2808 ? 1'h1 : _T_943;	// matmul/matmul-hw.mlir:8029:13, :13515:12, :17133:13
  assign _T_1863 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13516:12
  assign _T_1862 = _T_2808 ? A_reg_bank82_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9897:19, :12297:32, :13517:12
  assign _T_1861 = _T_2819 ? 1'h1 : _T_938;	// matmul/matmul-hw.mlir:8029:13, :13518:12, :17163:13
  assign _T_1860 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13519:12
  assign _T_1859 = _T_2819 ? A_reg_bank83_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9894:19, :12298:32, :13520:12
  assign _T_1858 = _T_2830 ? 1'h1 : _T_933;	// matmul/matmul-hw.mlir:8029:13, :13521:12, :17193:13
  assign _T_1857 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13522:12
  assign _T_1856 = _T_2830 ? A_reg_bank84_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9891:19, :12299:32, :13523:12
  assign _T_1855 = _T_2841 ? 1'h1 : _T_928;	// matmul/matmul-hw.mlir:8029:13, :13524:12, :17223:13
  assign _T_1854 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13525:12
  assign _T_1853 = _T_2841 ? A_reg_bank85_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9888:19, :12300:32, :13526:12
  assign _T_1852 = _T_2852 ? 1'h1 : _T_923;	// matmul/matmul-hw.mlir:8029:13, :13527:12, :17253:13
  assign _T_1851 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13528:12
  assign _T_1850 = _T_2852 ? A_reg_bank86_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9885:19, :12301:32, :13529:12
  assign _T_1849 = _T_2863 ? 1'h1 : _T_918;	// matmul/matmul-hw.mlir:8029:13, :13530:12, :17283:13
  assign _T_1848 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13531:12
  assign _T_1847 = _T_2863 ? A_reg_bank87_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9882:19, :12302:32, :13532:12
  assign _T_1846 = _T_2874 ? 1'h1 : _T_913;	// matmul/matmul-hw.mlir:8029:13, :13533:12, :17313:13
  assign _T_1845 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13534:12
  assign _T_1844 = _T_2874 ? A_reg_bank88_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9879:19, :12303:32, :13535:12
  assign _T_1843 = _T_2885 ? 1'h1 : _T_908;	// matmul/matmul-hw.mlir:8029:13, :13536:12, :17343:13
  assign _T_1842 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13537:12
  assign _T_1841 = _T_2885 ? A_reg_bank89_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9876:19, :12304:32, :13538:12
  assign _T_1840 = _T_2892 ? 1'h1 : _T_903;	// matmul/matmul-hw.mlir:8029:13, :13539:12, :17373:13
  assign _T_1839 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13540:12
  assign _T_1838 = _T_2892 ? A_reg_bank90_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9873:19, :12305:32, :13541:12
  assign _T_1837 = _T_2897 ? 1'h1 : _T_898;	// matmul/matmul-hw.mlir:8029:13, :13542:12, :17403:13
  assign _T_1836 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13543:12
  assign _T_1835 = _T_2897 ? A_reg_bank91_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9870:19, :12306:32, :13544:12
  assign _T_1834 = _T_2902 ? 1'h1 : _T_893;	// matmul/matmul-hw.mlir:8029:13, :13545:12, :17433:13
  assign _T_1833 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13546:12
  assign _T_1832 = _T_2902 ? A_reg_bank92_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9867:19, :12307:32, :13547:12
  assign _T_1831 = _T_2907 ? 1'h1 : _T_888;	// matmul/matmul-hw.mlir:8029:13, :13548:12, :17463:13
  assign _T_1830 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13549:12
  assign _T_1829 = _T_2907 ? A_reg_bank93_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9864:19, :12308:32, :13550:12
  assign _T_1828 = _T_2912 ? 1'h1 : _T_883;	// matmul/matmul-hw.mlir:8029:13, :13551:12, :17493:13
  assign _T_1827 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13552:12
  assign _T_1826 = _T_2912 ? A_reg_bank94_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9861:19, :12309:32, :13553:12
  wire [21:0] _T_2914 = _T_2913;	// matmul/matmul-hw.mlir:13555:12
  wire [21:0] _T_2915 = {_T_2914[5'h0+:21], {{_T_2712}}};	// matmul/matmul-hw.mlir:13556:19, :13557:12, :13558:12, :13559:12
  wire [21:0] _T_2916 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13560:19, :13561:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13562:5
    if (rst)	// matmul/matmul-hw.mlir:13562:5
      _T_2913 <= _T_2916;	// matmul/matmul-hw.mlir:13565:7
    else	// matmul/matmul-hw.mlir:13562:5
      _T_2913 <= _T_2915;	// matmul/matmul-hw.mlir:13563:7
  end // always @(posedge)
  wire _T_2917 = _T_2913[5'h15];	// matmul/matmul-hw.mlir:13555:12, :13567:16, :13568:12
  assign _T_1825 = _T_2917 ? 1'h1 : _T_878;	// matmul/matmul-hw.mlir:8029:13, :13569:12, :17523:13
  assign _T_1824 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13570:12
  assign _T_1823 = _T_2917 ? A_reg_bank95_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9858:19, :12310:32, :13571:12
  assign _T_1822 = _T_2797 ? 1'h1 : _T_866;	// matmul/matmul-hw.mlir:8029:13, :13572:12, :17668:13
  assign _T_1821 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13573:12
  assign _T_1820 = _T_2797 ? A_reg_bank96_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9855:19, :12311:32, :13574:12
  assign _T_1819 = _T_2808 ? 1'h1 : _T_861;	// matmul/matmul-hw.mlir:8029:13, :13575:12, :17698:13
  assign _T_1818 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13576:12
  assign _T_1817 = _T_2808 ? A_reg_bank97_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9852:19, :12312:32, :13577:12
  assign _T_1816 = _T_2819 ? 1'h1 : _T_856;	// matmul/matmul-hw.mlir:8029:13, :13578:12, :17728:13
  assign _T_1815 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13579:12
  assign _T_1814 = _T_2819 ? A_reg_bank98_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9849:19, :12313:32, :13580:12
  assign _T_1813 = _T_2830 ? 1'h1 : _T_851;	// matmul/matmul-hw.mlir:8029:13, :13581:12, :17758:13
  assign _T_1812 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13582:12
  assign _T_1811 = _T_2830 ? A_reg_bank99_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9846:19, :12314:32, :13583:12
  assign _T_1810 = _T_2841 ? 1'h1 : _T_846;	// matmul/matmul-hw.mlir:8029:13, :13584:12, :17788:13
  assign _T_1809 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13585:12
  assign _T_1808 = _T_2841 ? A_reg_bank100_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9843:19, :12315:33, :13586:12
  assign _T_1807 = _T_2852 ? 1'h1 : _T_841;	// matmul/matmul-hw.mlir:8029:13, :13587:12, :17818:13
  assign _T_1806 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13588:12
  assign _T_1805 = _T_2852 ? A_reg_bank101_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9840:19, :12316:33, :13589:12
  assign _T_1804 = _T_2863 ? 1'h1 : _T_836;	// matmul/matmul-hw.mlir:8029:13, :13590:12, :17848:13
  assign _T_1803 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13591:12
  assign _T_1802 = _T_2863 ? A_reg_bank102_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9837:19, :12317:33, :13592:12
  assign _T_1801 = _T_2874 ? 1'h1 : _T_831;	// matmul/matmul-hw.mlir:8029:13, :13593:12, :17878:13
  assign _T_1800 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13594:12
  assign _T_1799 = _T_2874 ? A_reg_bank103_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9834:19, :12318:33, :13595:12
  assign _T_1798 = _T_2885 ? 1'h1 : _T_826;	// matmul/matmul-hw.mlir:8029:13, :13596:12, :17908:13
  assign _T_1797 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13597:12
  assign _T_1796 = _T_2885 ? A_reg_bank104_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9831:19, :12319:33, :13598:12
  assign _T_1795 = _T_2892 ? 1'h1 : _T_821;	// matmul/matmul-hw.mlir:8029:13, :13599:12, :17938:13
  assign _T_1794 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13600:12
  assign _T_1793 = _T_2892 ? A_reg_bank105_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9828:19, :12320:33, :13601:12
  assign _T_1792 = _T_2897 ? 1'h1 : _T_816;	// matmul/matmul-hw.mlir:8029:13, :13602:12, :17968:13
  assign _T_1791 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13603:12
  assign _T_1790 = _T_2897 ? A_reg_bank106_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9825:19, :12321:33, :13604:12
  assign _T_1789 = _T_2902 ? 1'h1 : _T_811;	// matmul/matmul-hw.mlir:8029:13, :13605:12, :17998:13
  assign _T_1788 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13606:12
  assign _T_1787 = _T_2902 ? A_reg_bank107_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9822:19, :12322:33, :13607:12
  assign _T_1786 = _T_2907 ? 1'h1 : _T_806;	// matmul/matmul-hw.mlir:8029:13, :13608:12, :18028:13
  assign _T_1785 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13609:12
  assign _T_1784 = _T_2907 ? A_reg_bank108_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9819:19, :12323:33, :13610:12
  assign _T_1783 = _T_2912 ? 1'h1 : _T_801;	// matmul/matmul-hw.mlir:8029:13, :13611:12, :18058:13
  assign _T_1782 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13612:12
  assign _T_1781 = _T_2912 ? A_reg_bank109_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9816:19, :12324:33, :13613:12
  assign _T_1780 = _T_2917 ? 1'h1 : _T_796;	// matmul/matmul-hw.mlir:8029:13, :13614:12, :18088:13
  assign _T_1779 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13615:12
  assign _T_1778 = _T_2917 ? A_reg_bank110_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9813:19, :12325:33, :13616:12
  wire [22:0] _T_2919 = _T_2918;	// matmul/matmul-hw.mlir:13618:12
  wire [22:0] _T_2920 = {_T_2919[5'h0+:22], {{_T_2712}}};	// matmul/matmul-hw.mlir:13619:19, :13620:12, :13621:12, :13622:12
  wire [22:0] _T_2921 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13623:19, :13624:12
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13625:5
    if (rst)	// matmul/matmul-hw.mlir:13625:5
      _T_2918 <= _T_2921;	// matmul/matmul-hw.mlir:13628:7
    else	// matmul/matmul-hw.mlir:13625:5
      _T_2918 <= _T_2920;	// matmul/matmul-hw.mlir:13626:7
  end // always @(posedge)
  wire _T_2922 = _T_2918[5'h16];	// matmul/matmul-hw.mlir:13618:12, :13630:16, :13631:12
  assign _T_1777 = _T_2922 ? 1'h1 : _T_791;	// matmul/matmul-hw.mlir:8029:13, :13632:12, :18118:13
  assign _T_1776 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13633:12
  assign _T_1775 = _T_2922 ? A_reg_bank111_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9810:19, :12326:33, :13634:12
  assign _T_1774 = _T_2808 ? 1'h1 : _T_779;	// matmul/matmul-hw.mlir:8029:13, :13635:12, :18263:13
  assign _T_1773 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13636:13
  assign _T_1772 = _T_2808 ? A_reg_bank112_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9807:19, :12327:33, :13637:13
  assign _T_1771 = _T_2819 ? 1'h1 : _T_774;	// matmul/matmul-hw.mlir:8029:13, :13638:13, :18293:13
  assign _T_1770 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13639:13
  assign _T_1769 = _T_2819 ? A_reg_bank113_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9804:19, :12328:33, :13640:13
  assign _T_1768 = _T_2830 ? 1'h1 : _T_769;	// matmul/matmul-hw.mlir:8029:13, :13641:13, :18323:13
  assign _T_1767 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13642:13
  assign _T_1766 = _T_2830 ? A_reg_bank114_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9801:19, :12329:33, :13643:13
  assign _T_1765 = _T_2841 ? 1'h1 : _T_764;	// matmul/matmul-hw.mlir:8029:13, :13644:13, :18353:13
  assign _T_1764 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13645:13
  assign _T_1763 = _T_2841 ? A_reg_bank115_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9798:19, :12330:33, :13646:13
  assign _T_1762 = _T_2852 ? 1'h1 : _T_759;	// matmul/matmul-hw.mlir:8029:13, :13647:13, :18383:13
  assign _T_1761 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13648:13
  assign _T_1760 = _T_2852 ? A_reg_bank116_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9795:19, :12331:33, :13649:13
  assign _T_1759 = _T_2863 ? 1'h1 : _T_754;	// matmul/matmul-hw.mlir:8029:13, :13650:13, :18413:13
  assign _T_1758 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13651:13
  assign _T_1757 = _T_2863 ? A_reg_bank117_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9792:19, :12332:33, :13652:13
  assign _T_1756 = _T_2874 ? 1'h1 : _T_749;	// matmul/matmul-hw.mlir:8029:13, :13653:13, :18443:13
  assign _T_1755 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13654:13
  assign _T_1754 = _T_2874 ? A_reg_bank118_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9789:19, :12333:33, :13655:13
  assign _T_1753 = _T_2885 ? 1'h1 : _T_744;	// matmul/matmul-hw.mlir:8029:13, :13656:13, :18473:13
  assign _T_1752 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13657:13
  assign _T_1751 = _T_2885 ? A_reg_bank119_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9786:19, :12334:33, :13658:13
  assign _T_1750 = _T_2892 ? 1'h1 : _T_739;	// matmul/matmul-hw.mlir:8029:13, :13659:13, :18503:13
  assign _T_1749 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13660:13
  assign _T_1748 = _T_2892 ? A_reg_bank120_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9783:19, :12335:33, :13661:13
  assign _T_1747 = _T_2897 ? 1'h1 : _T_734;	// matmul/matmul-hw.mlir:8029:13, :13662:13, :18533:13
  assign _T_1746 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13663:13
  assign _T_1745 = _T_2897 ? A_reg_bank121_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9780:19, :12336:33, :13664:13
  assign _T_1744 = _T_2902 ? 1'h1 : _T_729;	// matmul/matmul-hw.mlir:8029:13, :13665:13, :18563:13
  assign _T_1743 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13666:13
  assign _T_1742 = _T_2902 ? A_reg_bank122_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9777:19, :12337:33, :13667:13
  assign _T_1741 = _T_2907 ? 1'h1 : _T_724;	// matmul/matmul-hw.mlir:8029:13, :13668:13, :18593:13
  assign _T_1740 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13669:13
  assign _T_1739 = _T_2907 ? A_reg_bank123_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9774:19, :12338:33, :13670:13
  assign _T_1738 = _T_2912 ? 1'h1 : _T_719;	// matmul/matmul-hw.mlir:8029:13, :13671:13, :18623:13
  assign _T_1737 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13672:13
  assign _T_1736 = _T_2912 ? A_reg_bank124_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9771:19, :12339:33, :13673:13
  assign _T_1735 = _T_2917 ? 1'h1 : _T_714;	// matmul/matmul-hw.mlir:8029:13, :13674:13, :18653:13
  assign _T_1734 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13675:13
  assign _T_1733 = _T_2917 ? A_reg_bank125_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9768:19, :12340:33, :13676:13
  assign _T_1732 = _T_2922 ? 1'h1 : _T_709;	// matmul/matmul-hw.mlir:8029:13, :13677:13, :18683:13
  assign _T_1731 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13678:13
  assign _T_1730 = _T_2922 ? A_reg_bank126_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9765:19, :12341:33, :13679:13
  wire [23:0] _T_2924 = _T_2923;	// matmul/matmul-hw.mlir:13681:13
  wire [23:0] _T_2925 = {_T_2924[5'h0+:23], {{_T_2712}}};	// matmul/matmul-hw.mlir:13682:19, :13683:13, :13684:13, :13685:13
  wire [23:0] _T_2926 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13686:19, :13687:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13688:5
    if (rst)	// matmul/matmul-hw.mlir:13688:5
      _T_2923 <= _T_2926;	// matmul/matmul-hw.mlir:13691:7
    else	// matmul/matmul-hw.mlir:13688:5
      _T_2923 <= _T_2925;	// matmul/matmul-hw.mlir:13689:7
  end // always @(posedge)
  wire _T_2927 = _T_2923[5'h17];	// matmul/matmul-hw.mlir:13681:13, :13693:15, :13694:13
  assign _T_1729 = _T_2927 ? 1'h1 : _T_704;	// matmul/matmul-hw.mlir:8029:13, :13695:13, :18713:13
  assign _T_1728 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13696:13
  assign _T_1727 = _T_2927 ? A_reg_bank127_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9762:19, :12342:33, :13697:13
  assign _T_1726 = _T_2819 ? 1'h1 : _T_692;	// matmul/matmul-hw.mlir:8029:13, :13698:13, :18858:13
  assign _T_1725 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13699:13
  assign _T_1724 = _T_2819 ? A_reg_bank128_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9759:19, :12343:33, :13700:13
  assign _T_1723 = _T_2830 ? 1'h1 : _T_687;	// matmul/matmul-hw.mlir:8029:13, :13701:13, :18888:13
  assign _T_1722 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13702:13
  assign _T_1721 = _T_2830 ? A_reg_bank129_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9756:19, :12344:33, :13703:13
  assign _T_1720 = _T_2841 ? 1'h1 : _T_682;	// matmul/matmul-hw.mlir:8029:13, :13704:13, :18918:13
  assign _T_1719 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13705:13
  assign _T_1718 = _T_2841 ? A_reg_bank130_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9753:19, :12345:33, :13706:13
  assign _T_1717 = _T_2852 ? 1'h1 : _T_677;	// matmul/matmul-hw.mlir:8029:13, :13707:13, :18948:13
  assign _T_1716 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13708:13
  assign _T_1715 = _T_2852 ? A_reg_bank131_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9750:19, :12346:33, :13709:13
  assign _T_1714 = _T_2863 ? 1'h1 : _T_672;	// matmul/matmul-hw.mlir:8029:13, :13710:13, :18978:13
  assign _T_1713 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13711:13
  assign _T_1712 = _T_2863 ? A_reg_bank132_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9747:19, :12347:33, :13712:13
  assign _T_1711 = _T_2874 ? 1'h1 : _T_667;	// matmul/matmul-hw.mlir:8029:13, :13713:13, :19008:13
  assign _T_1710 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13714:13
  assign _T_1709 = _T_2874 ? A_reg_bank133_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9744:19, :12348:33, :13715:13
  assign _T_1708 = _T_2885 ? 1'h1 : _T_662;	// matmul/matmul-hw.mlir:8029:13, :13716:13, :19038:13
  assign _T_1707 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13717:13
  assign _T_1706 = _T_2885 ? A_reg_bank134_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9741:19, :12349:33, :13718:13
  assign _T_1705 = _T_2892 ? 1'h1 : _T_657;	// matmul/matmul-hw.mlir:8029:13, :13719:13, :19068:13
  assign _T_1704 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13720:13
  assign _T_1703 = _T_2892 ? A_reg_bank135_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9738:19, :12350:33, :13721:13
  assign _T_1702 = _T_2897 ? 1'h1 : _T_652;	// matmul/matmul-hw.mlir:8029:13, :13722:13, :19098:13
  assign _T_1701 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13723:13
  assign _T_1700 = _T_2897 ? A_reg_bank136_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9735:19, :12351:33, :13724:13
  assign _T_1699 = _T_2902 ? 1'h1 : _T_647;	// matmul/matmul-hw.mlir:8029:13, :13725:13, :19128:13
  assign _T_1698 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13726:13
  assign _T_1697 = _T_2902 ? A_reg_bank137_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9732:19, :12352:33, :13727:13
  assign _T_1696 = _T_2907 ? 1'h1 : _T_642;	// matmul/matmul-hw.mlir:8029:13, :13728:13, :19158:13
  assign _T_1695 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13729:13
  assign _T_1694 = _T_2907 ? A_reg_bank138_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9729:19, :12353:33, :13730:13
  assign _T_1693 = _T_2912 ? 1'h1 : _T_637;	// matmul/matmul-hw.mlir:8029:13, :13731:13, :19188:13
  assign _T_1692 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13732:13
  assign _T_1691 = _T_2912 ? A_reg_bank139_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9726:19, :12354:33, :13733:13
  assign _T_1690 = _T_2917 ? 1'h1 : _T_632;	// matmul/matmul-hw.mlir:8029:13, :13734:13, :19218:13
  assign _T_1689 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13735:13
  assign _T_1688 = _T_2917 ? A_reg_bank140_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9723:19, :12355:33, :13736:13
  assign _T_1687 = _T_2922 ? 1'h1 : _T_627;	// matmul/matmul-hw.mlir:8029:13, :13737:13, :19248:13
  assign _T_1686 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13738:13
  assign _T_1685 = _T_2922 ? A_reg_bank141_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9720:19, :12356:33, :13739:13
  assign _T_1684 = _T_2927 ? 1'h1 : _T_622;	// matmul/matmul-hw.mlir:8029:13, :13740:13, :19278:13
  assign _T_1683 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13741:13
  assign _T_1682 = _T_2927 ? A_reg_bank142_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9717:19, :12357:33, :13742:13
  wire [24:0] _T_2929 = _T_2928;	// matmul/matmul-hw.mlir:13744:13
  wire [24:0] _T_2930 = {_T_2929[5'h0+:24], {{_T_2712}}};	// matmul/matmul-hw.mlir:13745:19, :13746:13, :13747:13, :13748:13
  wire [24:0] _T_2931 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13749:19, :13750:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13751:5
    if (rst)	// matmul/matmul-hw.mlir:13751:5
      _T_2928 <= _T_2931;	// matmul/matmul-hw.mlir:13754:7
    else	// matmul/matmul-hw.mlir:13751:5
      _T_2928 <= _T_2930;	// matmul/matmul-hw.mlir:13752:7
  end // always @(posedge)
  wire _T_2932 = _T_2928[5'h18];	// matmul/matmul-hw.mlir:13744:13, :13756:15, :13757:13
  assign _T_1681 = _T_2932 ? 1'h1 : _T_617;	// matmul/matmul-hw.mlir:8029:13, :13758:13, :19308:13
  assign _T_1680 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13759:13
  assign _T_1679 = _T_2932 ? A_reg_bank143_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9714:19, :12358:33, :13760:13
  assign _T_1678 = _T_2830 ? 1'h1 : _T_605;	// matmul/matmul-hw.mlir:8029:13, :13761:13, :19453:13
  assign _T_1677 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13762:13
  assign _T_1676 = _T_2830 ? A_reg_bank144_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9711:19, :12359:33, :13763:13
  assign _T_1675 = _T_2841 ? 1'h1 : _T_600;	// matmul/matmul-hw.mlir:8029:13, :13764:13, :19483:13
  assign _T_1674 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13765:13
  assign _T_1673 = _T_2841 ? A_reg_bank145_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9708:19, :12360:33, :13766:13
  assign _T_1672 = _T_2852 ? 1'h1 : _T_595;	// matmul/matmul-hw.mlir:8029:13, :13767:13, :19513:13
  assign _T_1671 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13768:13
  assign _T_1670 = _T_2852 ? A_reg_bank146_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9705:19, :12361:33, :13769:13
  assign _T_1669 = _T_2863 ? 1'h1 : _T_590;	// matmul/matmul-hw.mlir:8029:13, :13770:13, :19543:13
  assign _T_1668 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13771:13
  assign _T_1667 = _T_2863 ? A_reg_bank147_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9702:19, :12362:33, :13772:13
  assign _T_1666 = _T_2874 ? 1'h1 : _T_585;	// matmul/matmul-hw.mlir:8029:13, :13773:13, :19573:13
  assign _T_1665 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13774:13
  assign _T_1664 = _T_2874 ? A_reg_bank148_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9699:19, :12363:33, :13775:13
  assign _T_1663 = _T_2885 ? 1'h1 : _T_580;	// matmul/matmul-hw.mlir:8029:13, :13776:13, :19603:13
  assign _T_1662 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13777:13
  assign _T_1661 = _T_2885 ? A_reg_bank149_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9696:19, :12364:33, :13778:13
  assign _T_1660 = _T_2892 ? 1'h1 : _T_575;	// matmul/matmul-hw.mlir:8029:13, :13779:13, :19633:13
  assign _T_1659 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13780:13
  assign _T_1658 = _T_2892 ? A_reg_bank150_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9693:19, :12365:33, :13781:13
  assign _T_1657 = _T_2897 ? 1'h1 : _T_570;	// matmul/matmul-hw.mlir:8029:13, :13782:13, :19663:13
  assign _T_1656 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13783:13
  assign _T_1655 = _T_2897 ? A_reg_bank151_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9690:19, :12366:33, :13784:13
  assign _T_1654 = _T_2902 ? 1'h1 : _T_565;	// matmul/matmul-hw.mlir:8029:13, :13785:13, :19693:13
  assign _T_1653 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13786:13
  assign _T_1652 = _T_2902 ? A_reg_bank152_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9687:19, :12367:33, :13787:13
  assign _T_1651 = _T_2907 ? 1'h1 : _T_560;	// matmul/matmul-hw.mlir:8029:13, :13788:13, :19723:13
  assign _T_1650 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13789:13
  assign _T_1649 = _T_2907 ? A_reg_bank153_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9684:19, :12368:33, :13790:13
  assign _T_1648 = _T_2912 ? 1'h1 : _T_555;	// matmul/matmul-hw.mlir:8029:13, :13791:13, :19753:13
  assign _T_1647 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13792:13
  assign _T_1646 = _T_2912 ? A_reg_bank154_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9681:19, :12369:33, :13793:13
  assign _T_1645 = _T_2917 ? 1'h1 : _T_550;	// matmul/matmul-hw.mlir:8029:13, :13794:13, :19783:13
  assign _T_1644 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13795:13
  assign _T_1643 = _T_2917 ? A_reg_bank155_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9678:19, :12370:33, :13796:13
  assign _T_1642 = _T_2922 ? 1'h1 : _T_545;	// matmul/matmul-hw.mlir:8029:13, :13797:13, :19813:13
  assign _T_1641 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13798:13
  assign _T_1640 = _T_2922 ? A_reg_bank156_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9675:19, :12371:33, :13799:13
  assign _T_1639 = _T_2927 ? 1'h1 : _T_540;	// matmul/matmul-hw.mlir:8029:13, :13800:13, :19843:13
  assign _T_1638 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13801:13
  assign _T_1637 = _T_2927 ? A_reg_bank157_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9672:19, :12372:33, :13802:13
  assign _T_1636 = _T_2932 ? 1'h1 : _T_535;	// matmul/matmul-hw.mlir:8029:13, :13803:13, :19873:13
  assign _T_1635 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13804:13
  assign _T_1634 = _T_2932 ? A_reg_bank158_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9669:19, :12373:33, :13805:13
  wire [25:0] _T_2934 = _T_2933;	// matmul/matmul-hw.mlir:13807:13
  wire [25:0] _T_2935 = {_T_2934[5'h0+:25], {{_T_2712}}};	// matmul/matmul-hw.mlir:13808:19, :13809:13, :13810:13, :13811:13
  wire [25:0] _T_2936 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13812:19, :13813:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13814:5
    if (rst)	// matmul/matmul-hw.mlir:13814:5
      _T_2933 <= _T_2936;	// matmul/matmul-hw.mlir:13817:7
    else	// matmul/matmul-hw.mlir:13814:5
      _T_2933 <= _T_2935;	// matmul/matmul-hw.mlir:13815:7
  end // always @(posedge)
  wire _T_2937 = _T_2933[5'h19];	// matmul/matmul-hw.mlir:13807:13, :13819:15, :13820:13
  assign _T_1633 = _T_2937 ? 1'h1 : _T_530;	// matmul/matmul-hw.mlir:8029:13, :13821:13, :19903:13
  assign _T_1632 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13822:13
  assign _T_1631 = _T_2937 ? A_reg_bank159_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9666:19, :12374:33, :13823:13
  assign _T_1630 = _T_2841 ? 1'h1 : _T_518;	// matmul/matmul-hw.mlir:8029:13, :13824:13, :20048:13
  assign _T_1629 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13825:13
  assign _T_1628 = _T_2841 ? A_reg_bank160_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9663:19, :12375:33, :13826:13
  assign _T_1627 = _T_2852 ? 1'h1 : _T_513;	// matmul/matmul-hw.mlir:8029:13, :13827:13, :20078:13
  assign _T_1626 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13828:13
  assign _T_1625 = _T_2852 ? A_reg_bank161_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9660:19, :12376:33, :13829:13
  assign _T_1624 = _T_2863 ? 1'h1 : _T_508;	// matmul/matmul-hw.mlir:8029:13, :13830:13, :20108:13
  assign _T_1623 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13831:13
  assign _T_1622 = _T_2863 ? A_reg_bank162_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9657:19, :12377:33, :13832:13
  assign _T_1621 = _T_2874 ? 1'h1 : _T_503;	// matmul/matmul-hw.mlir:8029:13, :13833:13, :20138:13
  assign _T_1620 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13834:13
  assign _T_1619 = _T_2874 ? A_reg_bank163_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9654:19, :12378:33, :13835:13
  assign _T_1618 = _T_2885 ? 1'h1 : _T_498;	// matmul/matmul-hw.mlir:8029:13, :13836:13, :20168:13
  assign _T_1617 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13837:13
  assign _T_1616 = _T_2885 ? A_reg_bank164_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9651:19, :12379:33, :13838:13
  assign _T_1615 = _T_2892 ? 1'h1 : _T_493;	// matmul/matmul-hw.mlir:8029:13, :13839:13, :20198:13
  assign _T_1614 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13840:13
  assign _T_1613 = _T_2892 ? A_reg_bank165_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9648:19, :12380:33, :13841:13
  assign _T_1612 = _T_2897 ? 1'h1 : _T_488;	// matmul/matmul-hw.mlir:8029:13, :13842:13, :20228:13
  assign _T_1611 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13843:13
  assign _T_1610 = _T_2897 ? A_reg_bank166_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9645:19, :12381:33, :13844:13
  assign _T_1609 = _T_2902 ? 1'h1 : _T_483;	// matmul/matmul-hw.mlir:8029:13, :13845:13, :20258:13
  assign _T_1608 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13846:13
  assign _T_1607 = _T_2902 ? A_reg_bank167_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9642:19, :12382:33, :13847:13
  assign _T_1606 = _T_2907 ? 1'h1 : _T_478;	// matmul/matmul-hw.mlir:8029:13, :13848:13, :20288:13
  assign _T_1605 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13849:13
  assign _T_1604 = _T_2907 ? A_reg_bank168_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9639:19, :12383:33, :13850:13
  assign _T_1603 = _T_2912 ? 1'h1 : _T_473;	// matmul/matmul-hw.mlir:8029:13, :13851:13, :20318:13
  assign _T_1602 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13852:13
  assign _T_1601 = _T_2912 ? A_reg_bank169_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9636:19, :12384:33, :13853:13
  assign _T_1600 = _T_2917 ? 1'h1 : _T_468;	// matmul/matmul-hw.mlir:8029:13, :13854:13, :20348:13
  assign _T_1599 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13855:13
  assign _T_1598 = _T_2917 ? A_reg_bank170_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9633:19, :12385:33, :13856:13
  assign _T_1597 = _T_2922 ? 1'h1 : _T_463;	// matmul/matmul-hw.mlir:8029:13, :13857:13, :20378:13
  assign _T_1596 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13858:13
  assign _T_1595 = _T_2922 ? A_reg_bank171_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9630:19, :12386:33, :13859:13
  assign _T_1594 = _T_2927 ? 1'h1 : _T_458;	// matmul/matmul-hw.mlir:8029:13, :13860:13, :20408:13
  assign _T_1593 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13861:13
  assign _T_1592 = _T_2927 ? A_reg_bank172_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9627:19, :12387:33, :13862:13
  assign _T_1591 = _T_2932 ? 1'h1 : _T_453;	// matmul/matmul-hw.mlir:8029:13, :13863:13, :20438:13
  assign _T_1590 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13864:13
  assign _T_1589 = _T_2932 ? A_reg_bank173_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9624:19, :12388:33, :13865:13
  assign _T_1588 = _T_2937 ? 1'h1 : _T_448;	// matmul/matmul-hw.mlir:8029:13, :13866:13, :20468:13
  assign _T_1587 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13867:13
  assign _T_1586 = _T_2937 ? A_reg_bank174_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9621:19, :12389:33, :13868:13
  wire [26:0] _T_2939 = _T_2938;	// matmul/matmul-hw.mlir:13870:13
  wire [26:0] _T_2940 = {_T_2939[5'h0+:26], {{_T_2712}}};	// matmul/matmul-hw.mlir:13871:19, :13872:13, :13873:13, :13874:13
  wire [26:0] _T_2941 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13875:19, :13876:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13877:5
    if (rst)	// matmul/matmul-hw.mlir:13877:5
      _T_2938 <= _T_2941;	// matmul/matmul-hw.mlir:13880:7
    else	// matmul/matmul-hw.mlir:13877:5
      _T_2938 <= _T_2940;	// matmul/matmul-hw.mlir:13878:7
  end // always @(posedge)
  wire _T_2942 = _T_2938[5'h1A];	// matmul/matmul-hw.mlir:13870:13, :13882:15, :13883:13
  assign _T_1585 = _T_2942 ? 1'h1 : _T_443;	// matmul/matmul-hw.mlir:8029:13, :13884:13, :20498:13
  assign _T_1584 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13885:13
  assign _T_1583 = _T_2942 ? A_reg_bank175_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9618:19, :12390:33, :13886:13
  assign _T_1582 = _T_2852 ? 1'h1 : _T_431;	// matmul/matmul-hw.mlir:8029:13, :13887:13, :20643:13
  assign _T_1581 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13888:13
  assign _T_1580 = _T_2852 ? A_reg_bank176_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9615:19, :12391:33, :13889:13
  assign _T_1579 = _T_2863 ? 1'h1 : _T_426;	// matmul/matmul-hw.mlir:8029:13, :13890:13, :20673:13
  assign _T_1578 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13891:13
  assign _T_1577 = _T_2863 ? A_reg_bank177_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9612:19, :12392:33, :13892:13
  assign _T_1576 = _T_2874 ? 1'h1 : _T_421;	// matmul/matmul-hw.mlir:8029:13, :13893:13, :20703:13
  assign _T_1575 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13894:13
  assign _T_1574 = _T_2874 ? A_reg_bank178_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9609:19, :12393:33, :13895:13
  assign _T_1573 = _T_2885 ? 1'h1 : _T_416;	// matmul/matmul-hw.mlir:8029:13, :13896:13, :20733:13
  assign _T_1572 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13897:13
  assign _T_1571 = _T_2885 ? A_reg_bank179_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9606:19, :12394:33, :13898:13
  assign _T_1570 = _T_2892 ? 1'h1 : _T_411;	// matmul/matmul-hw.mlir:8029:13, :13899:13, :20763:13
  assign _T_1569 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13900:13
  assign _T_1568 = _T_2892 ? A_reg_bank180_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9603:19, :12395:33, :13901:13
  assign _T_1567 = _T_2897 ? 1'h1 : _T_406;	// matmul/matmul-hw.mlir:8029:13, :13902:13, :20793:13
  assign _T_1566 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13903:13
  assign _T_1565 = _T_2897 ? A_reg_bank181_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9600:19, :12396:33, :13904:13
  assign _T_1564 = _T_2902 ? 1'h1 : _T_401;	// matmul/matmul-hw.mlir:8029:13, :13905:13, :20823:13
  assign _T_1563 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13906:13
  assign _T_1562 = _T_2902 ? A_reg_bank182_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9597:19, :12397:33, :13907:13
  assign _T_1561 = _T_2907 ? 1'h1 : _T_396;	// matmul/matmul-hw.mlir:8029:13, :13908:13, :20853:13
  assign _T_1560 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13909:13
  assign _T_1559 = _T_2907 ? A_reg_bank183_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9594:19, :12398:33, :13910:13
  assign _T_1558 = _T_2912 ? 1'h1 : _T_391;	// matmul/matmul-hw.mlir:8029:13, :13911:13, :20883:13
  assign _T_1557 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13912:13
  assign _T_1556 = _T_2912 ? A_reg_bank184_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9591:19, :12399:33, :13913:13
  assign _T_1555 = _T_2917 ? 1'h1 : _T_386;	// matmul/matmul-hw.mlir:8029:13, :13914:13, :20913:13
  assign _T_1554 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13915:13
  assign _T_1553 = _T_2917 ? A_reg_bank185_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9588:19, :12400:33, :13916:13
  assign _T_1552 = _T_2922 ? 1'h1 : _T_381;	// matmul/matmul-hw.mlir:8029:13, :13917:13, :20943:13
  assign _T_1551 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13918:13
  assign _T_1550 = _T_2922 ? A_reg_bank186_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9585:19, :12401:33, :13919:13
  assign _T_1549 = _T_2927 ? 1'h1 : _T_376;	// matmul/matmul-hw.mlir:8029:13, :13920:13, :20973:13
  assign _T_1548 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13921:13
  assign _T_1547 = _T_2927 ? A_reg_bank187_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9582:19, :12402:33, :13922:13
  assign _T_1546 = _T_2932 ? 1'h1 : _T_371;	// matmul/matmul-hw.mlir:8029:13, :13923:13, :21003:13
  assign _T_1545 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13924:13
  assign _T_1544 = _T_2932 ? A_reg_bank188_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9579:19, :12403:33, :13925:13
  assign _T_1543 = _T_2937 ? 1'h1 : _T_366;	// matmul/matmul-hw.mlir:8029:13, :13926:13, :21033:13
  assign _T_1542 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13927:13
  assign _T_1541 = _T_2937 ? A_reg_bank189_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9576:19, :12404:33, :13928:13
  assign _T_1540 = _T_2942 ? 1'h1 : _T_361;	// matmul/matmul-hw.mlir:8029:13, :13929:13, :21063:13
  assign _T_1539 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13930:13
  assign _T_1538 = _T_2942 ? A_reg_bank190_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9573:19, :12405:33, :13931:13
  wire [27:0] _T_2944 = _T_2943;	// matmul/matmul-hw.mlir:13933:13
  wire [27:0] _T_2945 = {_T_2944[5'h0+:27], {{_T_2712}}};	// matmul/matmul-hw.mlir:13934:19, :13935:13, :13936:13, :13937:13
  wire [27:0] _T_2946 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:13938:19, :13939:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:13940:5
    if (rst)	// matmul/matmul-hw.mlir:13940:5
      _T_2943 <= _T_2946;	// matmul/matmul-hw.mlir:13943:7
    else	// matmul/matmul-hw.mlir:13940:5
      _T_2943 <= _T_2945;	// matmul/matmul-hw.mlir:13941:7
  end // always @(posedge)
  wire _T_2947 = _T_2943[5'h1B];	// matmul/matmul-hw.mlir:13933:13, :13945:15, :13946:13
  assign _T_1537 = _T_2947 ? 1'h1 : _T_356;	// matmul/matmul-hw.mlir:8029:13, :13947:13, :21093:13
  assign _T_1536 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13948:13
  assign _T_1535 = _T_2947 ? A_reg_bank191_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9570:19, :12406:33, :13949:13
  assign _T_1534 = _T_2863 ? 1'h1 : _T_344;	// matmul/matmul-hw.mlir:8029:13, :13950:13, :21238:13
  assign _T_1533 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13951:13
  assign _T_1532 = _T_2863 ? A_reg_bank192_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9567:19, :12407:33, :13952:13
  assign _T_1531 = _T_2874 ? 1'h1 : _T_339;	// matmul/matmul-hw.mlir:8029:13, :13953:13, :21268:13
  assign _T_1530 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13954:13
  assign _T_1529 = _T_2874 ? A_reg_bank193_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9564:19, :12408:33, :13955:13
  assign _T_1528 = _T_2885 ? 1'h1 : _T_334;	// matmul/matmul-hw.mlir:8029:13, :13956:13, :21298:13
  assign _T_1527 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13957:13
  assign _T_1526 = _T_2885 ? A_reg_bank194_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9561:19, :12409:33, :13958:13
  assign _T_1525 = _T_2892 ? 1'h1 : _T_329;	// matmul/matmul-hw.mlir:8029:13, :13959:13, :21328:13
  assign _T_1524 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13960:13
  assign _T_1523 = _T_2892 ? A_reg_bank195_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9558:19, :12410:33, :13961:13
  assign _T_1522 = _T_2897 ? 1'h1 : _T_324;	// matmul/matmul-hw.mlir:8029:13, :13962:13, :21358:13
  assign _T_1521 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13963:13
  assign _T_1520 = _T_2897 ? A_reg_bank196_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9555:19, :12411:33, :13964:13
  assign _T_1519 = _T_2902 ? 1'h1 : _T_319;	// matmul/matmul-hw.mlir:8029:13, :13965:13, :21388:13
  assign _T_1518 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13966:13
  assign _T_1517 = _T_2902 ? A_reg_bank197_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9552:19, :12412:33, :13967:13
  assign _T_1516 = _T_2907 ? 1'h1 : _T_314;	// matmul/matmul-hw.mlir:8029:13, :13968:13, :21418:13
  assign _T_1515 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13969:13
  assign _T_1514 = _T_2907 ? A_reg_bank198_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9549:19, :12413:33, :13970:13
  assign _T_1513 = _T_2912 ? 1'h1 : _T_309;	// matmul/matmul-hw.mlir:8029:13, :13971:13, :21448:13
  assign _T_1512 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13972:13
  assign _T_1511 = _T_2912 ? A_reg_bank199_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9546:19, :12414:33, :13973:13
  assign _T_1510 = _T_2917 ? 1'h1 : _T_304;	// matmul/matmul-hw.mlir:8029:13, :13974:13, :21478:13
  assign _T_1509 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13975:13
  assign _T_1508 = _T_2917 ? A_reg_bank200_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9543:19, :12415:33, :13976:13
  assign _T_1507 = _T_2922 ? 1'h1 : _T_299;	// matmul/matmul-hw.mlir:8029:13, :13977:13, :21508:13
  assign _T_1506 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13978:13
  assign _T_1505 = _T_2922 ? A_reg_bank201_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9540:19, :12416:33, :13979:13
  assign _T_1504 = _T_2927 ? 1'h1 : _T_294;	// matmul/matmul-hw.mlir:8029:13, :13980:13, :21538:13
  assign _T_1503 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13981:13
  assign _T_1502 = _T_2927 ? A_reg_bank202_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9537:19, :12417:33, :13982:13
  assign _T_1501 = _T_2932 ? 1'h1 : _T_289;	// matmul/matmul-hw.mlir:8029:13, :13983:13, :21568:13
  assign _T_1500 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13984:13
  assign _T_1499 = _T_2932 ? A_reg_bank203_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9534:19, :12418:33, :13985:13
  assign _T_1498 = _T_2937 ? 1'h1 : _T_284;	// matmul/matmul-hw.mlir:8029:13, :13986:13, :21598:13
  assign _T_1497 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13987:13
  assign _T_1496 = _T_2937 ? A_reg_bank204_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9531:19, :12419:33, :13988:13
  assign _T_1495 = _T_2942 ? 1'h1 : _T_279;	// matmul/matmul-hw.mlir:8029:13, :13989:13, :21628:13
  assign _T_1494 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13990:13
  assign _T_1493 = _T_2942 ? A_reg_bank205_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9528:19, :12420:33, :13991:13
  assign _T_1492 = _T_2947 ? 1'h1 : _T_274;	// matmul/matmul-hw.mlir:8029:13, :13992:13, :21658:13
  assign _T_1491 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :13993:13
  assign _T_1490 = _T_2947 ? A_reg_bank206_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9525:19, :12421:33, :13994:13
  wire [28:0] _T_2949 = _T_2948;	// matmul/matmul-hw.mlir:13996:13
  wire [28:0] _T_2950 = {_T_2949[5'h0+:28], {{_T_2712}}};	// matmul/matmul-hw.mlir:13997:19, :13998:13, :13999:13, :14000:13
  wire [28:0] _T_2951 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:14001:19, :14002:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14003:5
    if (rst)	// matmul/matmul-hw.mlir:14003:5
      _T_2948 <= _T_2951;	// matmul/matmul-hw.mlir:14006:7
    else	// matmul/matmul-hw.mlir:14003:5
      _T_2948 <= _T_2950;	// matmul/matmul-hw.mlir:14004:7
  end // always @(posedge)
  wire _T_2952 = _T_2948[5'h1C];	// matmul/matmul-hw.mlir:13996:13, :14008:15, :14009:13
  assign _T_1489 = _T_2952 ? 1'h1 : _T_269;	// matmul/matmul-hw.mlir:8029:13, :14010:13, :21688:13
  assign _T_1488 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14011:13
  assign _T_1487 = _T_2952 ? A_reg_bank207_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9522:19, :12422:33, :14012:13
  assign _T_1486 = _T_2874 ? 1'h1 : _T_257;	// matmul/matmul-hw.mlir:8029:13, :14013:13, :21848:13
  assign _T_1485 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14014:13
  assign _T_1484 = _T_2874 ? A_reg_bank208_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9519:19, :12423:33, :14015:13
  assign _T_1483 = _T_2885 ? 1'h1 : _T_252;	// matmul/matmul-hw.mlir:8029:13, :14016:13, :21878:13
  assign _T_1482 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14017:13
  assign _T_1481 = _T_2885 ? A_reg_bank209_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9516:19, :12424:33, :14018:13
  assign _T_1480 = _T_2892 ? 1'h1 : _T_247;	// matmul/matmul-hw.mlir:8029:13, :14019:13, :21908:13
  assign _T_1479 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14020:13
  assign _T_1478 = _T_2892 ? A_reg_bank210_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9513:19, :12425:33, :14021:13
  assign _T_1477 = _T_2897 ? 1'h1 : _T_242;	// matmul/matmul-hw.mlir:8029:13, :14022:13, :21938:13
  assign _T_1476 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14023:13
  assign _T_1475 = _T_2897 ? A_reg_bank211_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9510:19, :12426:33, :14024:13
  assign _T_1474 = _T_2902 ? 1'h1 : _T_237;	// matmul/matmul-hw.mlir:8029:13, :14025:13, :21968:13
  assign _T_1473 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14026:13
  assign _T_1472 = _T_2902 ? A_reg_bank212_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9507:19, :12427:33, :14027:13
  assign _T_1471 = _T_2907 ? 1'h1 : _T_232;	// matmul/matmul-hw.mlir:8029:13, :14028:13, :21998:13
  assign _T_1470 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14029:13
  assign _T_1469 = _T_2907 ? A_reg_bank213_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9504:19, :12428:33, :14030:13
  assign _T_1468 = _T_2912 ? 1'h1 : _T_227;	// matmul/matmul-hw.mlir:8029:13, :14031:13, :22028:13
  assign _T_1467 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14032:13
  assign _T_1466 = _T_2912 ? A_reg_bank214_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9501:19, :12429:33, :14033:13
  assign _T_1465 = _T_2917 ? 1'h1 : _T_222;	// matmul/matmul-hw.mlir:8029:13, :14034:13, :22058:13
  assign _T_1464 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14035:13
  assign _T_1463 = _T_2917 ? A_reg_bank215_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9498:19, :12430:33, :14036:13
  assign _T_1462 = _T_2922 ? 1'h1 : _T_217;	// matmul/matmul-hw.mlir:8029:13, :14037:13, :22088:13
  assign _T_1461 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14038:13
  assign _T_1460 = _T_2922 ? A_reg_bank216_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9495:19, :12431:33, :14039:13
  assign _T_1459 = _T_2927 ? 1'h1 : _T_212;	// matmul/matmul-hw.mlir:8029:13, :14040:13, :22118:13
  assign _T_1458 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14041:13
  assign _T_1457 = _T_2927 ? A_reg_bank217_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9492:19, :12432:33, :14042:13
  assign _T_1456 = _T_2932 ? 1'h1 : _T_207;	// matmul/matmul-hw.mlir:8029:13, :14043:13, :22148:13
  assign _T_1455 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14044:13
  assign _T_1454 = _T_2932 ? A_reg_bank218_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9489:19, :12433:33, :14045:13
  assign _T_1453 = _T_2937 ? 1'h1 : _T_202;	// matmul/matmul-hw.mlir:8029:13, :14046:13, :22178:13
  assign _T_1452 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14047:13
  assign _T_1451 = _T_2937 ? A_reg_bank219_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9486:19, :12434:33, :14048:13
  assign _T_1450 = _T_2942 ? 1'h1 : _T_197;	// matmul/matmul-hw.mlir:8029:13, :14049:13, :22208:13
  assign _T_1449 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14050:13
  assign _T_1448 = _T_2942 ? A_reg_bank220_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9483:19, :12435:33, :14051:13
  assign _T_1447 = _T_2947 ? 1'h1 : _T_192;	// matmul/matmul-hw.mlir:8029:13, :14052:13, :22238:13
  assign _T_1446 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14053:13
  assign _T_1445 = _T_2947 ? A_reg_bank221_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9480:19, :12436:33, :14054:13
  assign _T_1444 = _T_2952 ? 1'h1 : _T_187;	// matmul/matmul-hw.mlir:8029:13, :14055:13, :22268:13
  assign _T_1443 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14056:13
  assign _T_1442 = _T_2952 ? A_reg_bank222_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9477:19, :12437:33, :14057:13
  wire [29:0] _T_2954 = _T_2953;	// matmul/matmul-hw.mlir:14059:13
  wire [29:0] _T_2955 = {_T_2954[5'h0+:29], {{_T_2712}}};	// matmul/matmul-hw.mlir:14060:19, :14061:13, :14062:13, :14063:13
  wire [29:0] _T_2956 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:14064:19, :14065:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14066:5
    if (rst)	// matmul/matmul-hw.mlir:14066:5
      _T_2953 <= _T_2956;	// matmul/matmul-hw.mlir:14069:7
    else	// matmul/matmul-hw.mlir:14066:5
      _T_2953 <= _T_2955;	// matmul/matmul-hw.mlir:14067:7
  end // always @(posedge)
  wire _T_2957 = _T_2953[5'h1D];	// matmul/matmul-hw.mlir:14059:13, :14071:15, :14072:13
  assign _T_1441 = _T_2957 ? 1'h1 : _T_182;	// matmul/matmul-hw.mlir:8029:13, :14073:13, :22298:13
  assign _T_1440 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14074:13
  assign _T_1439 = _T_2957 ? A_reg_bank223_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9474:19, :12438:33, :14075:13
  assign _T_1438 = _T_2885 ? 1'h1 : _T_170;	// matmul/matmul-hw.mlir:8029:13, :14076:13, :22458:13
  assign _T_1437 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14077:13
  assign _T_1436 = _T_2885 ? A_reg_bank224_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9471:19, :12439:33, :14078:13
  assign _T_1435 = _T_2892 ? 1'h1 : _T_165;	// matmul/matmul-hw.mlir:8029:13, :14079:13, :22488:13
  assign _T_1434 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14080:13
  assign _T_1433 = _T_2892 ? A_reg_bank225_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9468:19, :12440:33, :14081:13
  assign _T_1432 = _T_2897 ? 1'h1 : _T_160;	// matmul/matmul-hw.mlir:8029:13, :14082:13, :22518:13
  assign _T_1431 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14083:13
  assign _T_1430 = _T_2897 ? A_reg_bank226_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9465:19, :12441:33, :14084:13
  assign _T_1429 = _T_2902 ? 1'h1 : _T_155;	// matmul/matmul-hw.mlir:8029:13, :14085:13, :22548:13
  assign _T_1428 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14086:13
  assign _T_1427 = _T_2902 ? A_reg_bank227_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9462:19, :12442:33, :14087:13
  assign _T_1426 = _T_2907 ? 1'h1 : _T_150;	// matmul/matmul-hw.mlir:8029:13, :14088:13, :22578:13
  assign _T_1425 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14089:13
  assign _T_1424 = _T_2907 ? A_reg_bank228_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9459:19, :12443:33, :14090:13
  assign _T_1423 = _T_2912 ? 1'h1 : _T_145;	// matmul/matmul-hw.mlir:8029:13, :14091:13, :22608:13
  assign _T_1422 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14092:13
  assign _T_1421 = _T_2912 ? A_reg_bank229_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9456:19, :12444:33, :14093:13
  assign _T_1420 = _T_2917 ? 1'h1 : _T_140;	// matmul/matmul-hw.mlir:8029:13, :14094:13, :22638:13
  assign _T_1419 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14095:13
  assign _T_1418 = _T_2917 ? A_reg_bank230_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9453:19, :12445:33, :14096:13
  assign _T_1417 = _T_2922 ? 1'h1 : _T_135;	// matmul/matmul-hw.mlir:8029:13, :14097:13, :22668:13
  assign _T_1416 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14098:13
  assign _T_1415 = _T_2922 ? A_reg_bank231_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9450:19, :12446:33, :14099:13
  assign _T_1414 = _T_2927 ? 1'h1 : _T_130;	// matmul/matmul-hw.mlir:8029:13, :14100:13, :22698:13
  assign _T_1413 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14101:13
  assign _T_1412 = _T_2927 ? A_reg_bank232_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9447:19, :12447:33, :14102:13
  assign _T_1411 = _T_2932 ? 1'h1 : _T_125;	// matmul/matmul-hw.mlir:8029:13, :14103:13, :22728:13
  assign _T_1410 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14104:13
  assign _T_1409 = _T_2932 ? A_reg_bank233_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9444:19, :12448:33, :14105:13
  assign _T_1408 = _T_2937 ? 1'h1 : _T_120;	// matmul/matmul-hw.mlir:8029:13, :14106:13, :22758:13
  assign _T_1407 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14107:13
  assign _T_1406 = _T_2937 ? A_reg_bank234_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9441:19, :12449:33, :14108:13
  assign _T_1405 = _T_2942 ? 1'h1 : _T_115;	// matmul/matmul-hw.mlir:8029:13, :14109:13, :22788:13
  assign _T_1404 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14110:13
  assign _T_1403 = _T_2942 ? A_reg_bank235_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9438:19, :12450:33, :14111:13
  assign _T_1402 = _T_2947 ? 1'h1 : _T_110;	// matmul/matmul-hw.mlir:8029:13, :14112:13, :22818:13
  assign _T_1401 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14113:13
  assign _T_1400 = _T_2947 ? A_reg_bank236_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9435:19, :12451:33, :14114:13
  assign _T_1399 = _T_2952 ? 1'h1 : _T_105;	// matmul/matmul-hw.mlir:8029:13, :14115:13, :22848:13
  assign _T_1398 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14116:13
  assign _T_1397 = _T_2952 ? A_reg_bank237_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9432:19, :12452:33, :14117:13
  assign _T_1396 = _T_2957 ? 1'h1 : _T_100;	// matmul/matmul-hw.mlir:8029:13, :14118:13, :22878:13
  assign _T_1395 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14119:13
  assign _T_1394 = _T_2957 ? A_reg_bank238_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9429:19, :12453:33, :14120:13
  wire [30:0] _T_2959 = _T_2958;	// matmul/matmul-hw.mlir:14122:13
  wire [30:0] _T_2960 = {_T_2959[5'h0+:30], {{_T_2712}}};	// matmul/matmul-hw.mlir:14123:19, :14124:13, :14125:13, :14126:13
  wire [30:0] _T_2961 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:14127:19, :14128:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14129:5
    if (rst)	// matmul/matmul-hw.mlir:14129:5
      _T_2958 <= _T_2961;	// matmul/matmul-hw.mlir:14132:7
    else	// matmul/matmul-hw.mlir:14129:5
      _T_2958 <= _T_2960;	// matmul/matmul-hw.mlir:14130:7
  end // always @(posedge)
  wire _T_2962 = _T_2958[5'h1E];	// matmul/matmul-hw.mlir:14122:13, :14134:15, :14135:13
  assign _T_1393 = _T_2962 ? 1'h1 : _T_95;	// matmul/matmul-hw.mlir:8029:13, :14136:13, :22908:13
  assign _T_1392 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14137:13
  assign _T_1391 = _T_2962 ? A_reg_bank239_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:9426:19, :12454:33, :14138:13
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0 (	// matmul/matmul-hw.mlir:14207:31
    .p0_rd_en   (_T_1386),	// matmul/matmul-hw.mlir:14229:13
    .p1_wr_en   (_T_1390),	// matmul/matmul-hw.mlir:14224:13
    .p1_wr_data (_T_1389),	// matmul/matmul-hw.mlir:14225:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2453)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1 (	// matmul/matmul-hw.mlir:14208:31
    .p0_rd_en   (_T_1381),	// matmul/matmul-hw.mlir:14251:13
    .p1_wr_en   (_T_1385),	// matmul/matmul-hw.mlir:14246:13
    .p1_wr_data (_T_1384),	// matmul/matmul-hw.mlir:14247:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2452)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2 (	// matmul/matmul-hw.mlir:14209:31
    .p0_rd_en   (_T_1376),	// matmul/matmul-hw.mlir:14273:13
    .p1_wr_en   (_T_1380),	// matmul/matmul-hw.mlir:14268:13
    .p1_wr_data (_T_1379),	// matmul/matmul-hw.mlir:14269:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2451)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3 (	// matmul/matmul-hw.mlir:14210:31
    .p0_rd_en   (_T_1371),	// matmul/matmul-hw.mlir:14295:13
    .p1_wr_en   (_T_1375),	// matmul/matmul-hw.mlir:14290:13
    .p1_wr_data (_T_1374),	// matmul/matmul-hw.mlir:14291:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2450)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4 (	// matmul/matmul-hw.mlir:14211:31
    .p0_rd_en   (_T_1366),	// matmul/matmul-hw.mlir:14317:13
    .p1_wr_en   (_T_1370),	// matmul/matmul-hw.mlir:14312:13
    .p1_wr_data (_T_1369),	// matmul/matmul-hw.mlir:14313:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2449)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5 (	// matmul/matmul-hw.mlir:14212:31
    .p0_rd_en   (_T_1361),	// matmul/matmul-hw.mlir:14339:13
    .p1_wr_en   (_T_1365),	// matmul/matmul-hw.mlir:14334:13
    .p1_wr_data (_T_1364),	// matmul/matmul-hw.mlir:14335:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2448)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6 (	// matmul/matmul-hw.mlir:14213:31
    .p0_rd_en   (_T_1356),	// matmul/matmul-hw.mlir:14361:13
    .p1_wr_en   (_T_1360),	// matmul/matmul-hw.mlir:14356:13
    .p1_wr_data (_T_1359),	// matmul/matmul-hw.mlir:14357:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2447)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7 (	// matmul/matmul-hw.mlir:14214:31
    .p0_rd_en   (_T_1351),	// matmul/matmul-hw.mlir:14383:13
    .p1_wr_en   (_T_1355),	// matmul/matmul-hw.mlir:14378:13
    .p1_wr_data (_T_1354),	// matmul/matmul-hw.mlir:14379:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2446)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8 (	// matmul/matmul-hw.mlir:14215:31
    .p0_rd_en   (_T_1346),	// matmul/matmul-hw.mlir:14405:13
    .p1_wr_en   (_T_1350),	// matmul/matmul-hw.mlir:14400:13
    .p1_wr_data (_T_1349),	// matmul/matmul-hw.mlir:14401:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2445)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9 (	// matmul/matmul-hw.mlir:14216:31
    .p0_rd_en   (_T_1341),	// matmul/matmul-hw.mlir:14427:13
    .p1_wr_en   (_T_1345),	// matmul/matmul-hw.mlir:14422:13
    .p1_wr_data (_T_1344),	// matmul/matmul-hw.mlir:14423:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2444)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10 (	// matmul/matmul-hw.mlir:14217:32
    .p0_rd_en   (_T_1336),	// matmul/matmul-hw.mlir:14449:13
    .p1_wr_en   (_T_1340),	// matmul/matmul-hw.mlir:14444:13
    .p1_wr_data (_T_1339),	// matmul/matmul-hw.mlir:14445:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2443)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11 (	// matmul/matmul-hw.mlir:14218:32
    .p0_rd_en   (_T_1331),	// matmul/matmul-hw.mlir:14471:13
    .p1_wr_en   (_T_1335),	// matmul/matmul-hw.mlir:14466:13
    .p1_wr_data (_T_1334),	// matmul/matmul-hw.mlir:14467:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2442)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12 (	// matmul/matmul-hw.mlir:14219:32
    .p0_rd_en   (_T_1326),	// matmul/matmul-hw.mlir:14493:13
    .p1_wr_en   (_T_1330),	// matmul/matmul-hw.mlir:14488:13
    .p1_wr_data (_T_1329),	// matmul/matmul-hw.mlir:14489:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2441)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13 (	// matmul/matmul-hw.mlir:14220:32
    .p0_rd_en   (_T_1321),	// matmul/matmul-hw.mlir:14515:13
    .p1_wr_en   (_T_1325),	// matmul/matmul-hw.mlir:14510:13
    .p1_wr_data (_T_1324),	// matmul/matmul-hw.mlir:14511:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2440)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14 (	// matmul/matmul-hw.mlir:14221:32
    .p0_rd_en   (_T_1316),	// matmul/matmul-hw.mlir:14537:13
    .p1_wr_en   (_T_1320),	// matmul/matmul-hw.mlir:14532:13
    .p1_wr_data (_T_1319),	// matmul/matmul-hw.mlir:14533:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2439)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15 (	// matmul/matmul-hw.mlir:14222:32
    .p0_rd_en   (_T_1311),	// matmul/matmul-hw.mlir:14559:13
    .p1_wr_en   (_T_1315),	// matmul/matmul-hw.mlir:14554:13
    .p1_wr_data (_T_1314),	// matmul/matmul-hw.mlir:14555:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2438)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16 (	// matmul/matmul-hw.mlir:14223:32
    .p0_rd_en   (_T_1308),	// matmul/matmul-hw.mlir:14578:13
    .p1_wr_en   (_T_1310),	// matmul/matmul-hw.mlir:14576:13
    .p1_wr_data (_T_1309),	// matmul/matmul-hw.mlir:14577:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2437)
  );
  assign _T_1390 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14224:13
  assign _T_1389 = _T_2742 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :9424:19, :14225:13
  assign _T_1388 = _T_2731 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14226:13
  assign _T_1387 = _T_2731 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14227:13
  mult mult_inst0 (	// matmul/matmul-hw.mlir:14228:26
    .a      (A_reg_bank0_p0_rd_data),	// matmul/matmul-hw.mlir:12215:31
    .b      (_T_2454),
    .t      (_T_2731),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst0_result)
  );
  assign _T_1386 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14229:13
  assign a_i_k_0_i_j_0 = A_reg_bank0_p0_rd_data;	// matmul/matmul-hw.mlir:12215:31, :14231:5
  //PROBE: a_i_k_0_i_j_0	// matmul/matmul-hw.mlir:14232:5
  assign b_i_k_0_i_j_0 = _T_2454;	// matmul/matmul-hw.mlir:14234:5
  //PROBE: b_i_k_0_i_j_0	// matmul/matmul-hw.mlir:14235:5
  assign c_prev_i_k_0_i_j_0 = C_reg_bank0_p0_rd_data_2453;	// matmul/matmul-hw.mlir:14207:31, :14237:5
  //PROBE: c_prev_i_k_0_i_j_0	// matmul/matmul-hw.mlir:14238:5
  assign tk_i_k_0_i_j_0 = _T_2712;	// matmul/matmul-hw.mlir:14240:5
  //PROBE: tk_i_k_0_i_j_0	// matmul/matmul-hw.mlir:14241:5
  wire [31:0] _T_2963 = mult_inst0_result + C_reg_bank0_p0_rd_data_2453;	// matmul/matmul-hw.mlir:14207:31, :14228:26, :14242:13
  assign c_i_k_0_i_j_0 = _T_2963;	// matmul/matmul-hw.mlir:14244:5
  //PROBE: c_i_k_0_i_j_0	// matmul/matmul-hw.mlir:14245:5
  assign _T_1385 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14246:13
  assign _T_1384 = _T_2753 ? _T_2963 : 32'bx;	// matmul/matmul-hw.mlir:9419:19, :14247:13
  assign _T_1383 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14248:13
  assign _T_1382 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14249:13
  mult mult_inst1 (	// matmul/matmul-hw.mlir:14250:26
    .a      (A_reg_bank1_p0_rd_data),	// matmul/matmul-hw.mlir:12216:31
    .b      (_T_2470),
    .t      (_T_2742),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst1_result)
  );
  assign _T_1381 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14251:13
  assign a_i_k_1_i_j_0 = A_reg_bank1_p0_rd_data;	// matmul/matmul-hw.mlir:12216:31, :14253:5
  //PROBE: a_i_k_1_i_j_0	// matmul/matmul-hw.mlir:14254:5
  assign b_i_k_1_i_j_0 = _T_2470;	// matmul/matmul-hw.mlir:14256:5
  //PROBE: b_i_k_1_i_j_0	// matmul/matmul-hw.mlir:14257:5
  assign c_prev_i_k_1_i_j_0 = C_reg_bank1_p0_rd_data_2452;	// matmul/matmul-hw.mlir:14208:31, :14259:5
  //PROBE: c_prev_i_k_1_i_j_0	// matmul/matmul-hw.mlir:14260:5
  assign tk_i_k_1_i_j_0 = _T_2189;	// matmul/matmul-hw.mlir:12484:12, :14262:5
  //PROBE: tk_i_k_1_i_j_0	// matmul/matmul-hw.mlir:14263:5
  wire [31:0] _T_2964 = mult_inst1_result + C_reg_bank1_p0_rd_data_2452;	// matmul/matmul-hw.mlir:14208:31, :14250:26, :14264:13
  assign c_i_k_1_i_j_0 = _T_2964;	// matmul/matmul-hw.mlir:14266:5
  //PROBE: c_i_k_1_i_j_0	// matmul/matmul-hw.mlir:14267:5
  assign _T_1380 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14268:13
  assign _T_1379 = _T_2764 ? _T_2964 : 32'bx;	// matmul/matmul-hw.mlir:9414:19, :14269:13
  assign _T_1378 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14270:13
  assign _T_1377 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14271:13
  mult mult_inst2 (	// matmul/matmul-hw.mlir:14272:26
    .a      (A_reg_bank2_p0_rd_data),	// matmul/matmul-hw.mlir:12217:31
    .b      (_T_2486),
    .t      (_T_2753),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst2_result)
  );
  assign _T_1376 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14273:13
  assign a_i_k_2_i_j_0 = A_reg_bank2_p0_rd_data;	// matmul/matmul-hw.mlir:12217:31, :14275:5
  //PROBE: a_i_k_2_i_j_0	// matmul/matmul-hw.mlir:14276:5
  assign b_i_k_2_i_j_0 = _T_2486;	// matmul/matmul-hw.mlir:14278:5
  //PROBE: b_i_k_2_i_j_0	// matmul/matmul-hw.mlir:14279:5
  assign c_prev_i_k_2_i_j_0 = C_reg_bank2_p0_rd_data_2451;	// matmul/matmul-hw.mlir:14209:31, :14281:5
  //PROBE: c_prev_i_k_2_i_j_0	// matmul/matmul-hw.mlir:14282:5
  assign tk_i_k_2_i_j_0 = _T_2731;	// matmul/matmul-hw.mlir:14284:5
  //PROBE: tk_i_k_2_i_j_0	// matmul/matmul-hw.mlir:14285:5
  wire [31:0] _T_2965 = mult_inst2_result + C_reg_bank2_p0_rd_data_2451;	// matmul/matmul-hw.mlir:14209:31, :14272:26, :14286:13
  assign c_i_k_2_i_j_0 = _T_2965;	// matmul/matmul-hw.mlir:14288:5
  //PROBE: c_i_k_2_i_j_0	// matmul/matmul-hw.mlir:14289:5
  assign _T_1375 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14290:13
  assign _T_1374 = _T_2775 ? _T_2965 : 32'bx;	// matmul/matmul-hw.mlir:9409:19, :14291:13
  assign _T_1373 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14292:13
  assign _T_1372 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14293:13
  mult mult_inst3 (	// matmul/matmul-hw.mlir:14294:26
    .a      (A_reg_bank3_p0_rd_data),	// matmul/matmul-hw.mlir:12218:31
    .b      (_T_2502),
    .t      (_T_2764),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst3_result)
  );
  assign _T_1371 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14295:13
  assign a_i_k_3_i_j_0 = A_reg_bank3_p0_rd_data;	// matmul/matmul-hw.mlir:12218:31, :14297:5
  //PROBE: a_i_k_3_i_j_0	// matmul/matmul-hw.mlir:14298:5
  assign b_i_k_3_i_j_0 = _T_2502;	// matmul/matmul-hw.mlir:14300:5
  //PROBE: b_i_k_3_i_j_0	// matmul/matmul-hw.mlir:14301:5
  assign c_prev_i_k_3_i_j_0 = C_reg_bank3_p0_rd_data_2450;	// matmul/matmul-hw.mlir:14210:31, :14303:5
  //PROBE: c_prev_i_k_3_i_j_0	// matmul/matmul-hw.mlir:14304:5
  assign tk_i_k_3_i_j_0 = _T_2742;	// matmul/matmul-hw.mlir:14306:5
  //PROBE: tk_i_k_3_i_j_0	// matmul/matmul-hw.mlir:14307:5
  wire [31:0] _T_2966 = mult_inst3_result + C_reg_bank3_p0_rd_data_2450;	// matmul/matmul-hw.mlir:14210:31, :14294:26, :14308:13
  assign c_i_k_3_i_j_0 = _T_2966;	// matmul/matmul-hw.mlir:14310:5
  //PROBE: c_i_k_3_i_j_0	// matmul/matmul-hw.mlir:14311:5
  assign _T_1370 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14312:13
  assign _T_1369 = _T_2786 ? _T_2966 : 32'bx;	// matmul/matmul-hw.mlir:9404:19, :14313:13
  assign _T_1368 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14314:13
  assign _T_1367 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14315:13
  mult mult_inst4 (	// matmul/matmul-hw.mlir:14316:26
    .a      (A_reg_bank4_p0_rd_data),	// matmul/matmul-hw.mlir:12219:31
    .b      (_T_2518),
    .t      (_T_2775),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst4_result)
  );
  assign _T_1366 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14317:13
  assign a_i_k_4_i_j_0 = A_reg_bank4_p0_rd_data;	// matmul/matmul-hw.mlir:12219:31, :14319:5
  //PROBE: a_i_k_4_i_j_0	// matmul/matmul-hw.mlir:14320:5
  assign b_i_k_4_i_j_0 = _T_2518;	// matmul/matmul-hw.mlir:14322:5
  //PROBE: b_i_k_4_i_j_0	// matmul/matmul-hw.mlir:14323:5
  assign c_prev_i_k_4_i_j_0 = C_reg_bank4_p0_rd_data_2449;	// matmul/matmul-hw.mlir:14211:31, :14325:5
  //PROBE: c_prev_i_k_4_i_j_0	// matmul/matmul-hw.mlir:14326:5
  assign tk_i_k_4_i_j_0 = _T_2753;	// matmul/matmul-hw.mlir:14328:5
  //PROBE: tk_i_k_4_i_j_0	// matmul/matmul-hw.mlir:14329:5
  wire [31:0] _T_2967 = mult_inst4_result + C_reg_bank4_p0_rd_data_2449;	// matmul/matmul-hw.mlir:14211:31, :14316:26, :14330:13
  assign c_i_k_4_i_j_0 = _T_2967;	// matmul/matmul-hw.mlir:14332:5
  //PROBE: c_i_k_4_i_j_0	// matmul/matmul-hw.mlir:14333:5
  assign _T_1365 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14334:13
  assign _T_1364 = _T_2797 ? _T_2967 : 32'bx;	// matmul/matmul-hw.mlir:9399:19, :14335:13
  assign _T_1363 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14336:13
  assign _T_1362 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14337:13
  mult mult_inst5 (	// matmul/matmul-hw.mlir:14338:26
    .a      (A_reg_bank5_p0_rd_data),	// matmul/matmul-hw.mlir:12220:31
    .b      (_T_2534),
    .t      (_T_2786),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst5_result)
  );
  assign _T_1361 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14339:13
  assign a_i_k_5_i_j_0 = A_reg_bank5_p0_rd_data;	// matmul/matmul-hw.mlir:12220:31, :14341:5
  //PROBE: a_i_k_5_i_j_0	// matmul/matmul-hw.mlir:14342:5
  assign b_i_k_5_i_j_0 = _T_2534;	// matmul/matmul-hw.mlir:14344:5
  //PROBE: b_i_k_5_i_j_0	// matmul/matmul-hw.mlir:14345:5
  assign c_prev_i_k_5_i_j_0 = C_reg_bank5_p0_rd_data_2448;	// matmul/matmul-hw.mlir:14212:31, :14347:5
  //PROBE: c_prev_i_k_5_i_j_0	// matmul/matmul-hw.mlir:14348:5
  assign tk_i_k_5_i_j_0 = _T_2764;	// matmul/matmul-hw.mlir:14350:5
  //PROBE: tk_i_k_5_i_j_0	// matmul/matmul-hw.mlir:14351:5
  wire [31:0] _T_2968 = mult_inst5_result + C_reg_bank5_p0_rd_data_2448;	// matmul/matmul-hw.mlir:14212:31, :14338:26, :14352:13
  assign c_i_k_5_i_j_0 = _T_2968;	// matmul/matmul-hw.mlir:14354:5
  //PROBE: c_i_k_5_i_j_0	// matmul/matmul-hw.mlir:14355:5
  assign _T_1360 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14356:13
  assign _T_1359 = _T_2808 ? _T_2968 : 32'bx;	// matmul/matmul-hw.mlir:9394:19, :14357:13
  assign _T_1358 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14358:13
  assign _T_1357 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14359:13
  mult mult_inst6 (	// matmul/matmul-hw.mlir:14360:26
    .a      (A_reg_bank6_p0_rd_data),	// matmul/matmul-hw.mlir:12221:31
    .b      (_T_2550),
    .t      (_T_2797),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst6_result)
  );
  assign _T_1356 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14361:13
  assign a_i_k_6_i_j_0 = A_reg_bank6_p0_rd_data;	// matmul/matmul-hw.mlir:12221:31, :14363:5
  //PROBE: a_i_k_6_i_j_0	// matmul/matmul-hw.mlir:14364:5
  assign b_i_k_6_i_j_0 = _T_2550;	// matmul/matmul-hw.mlir:14366:5
  //PROBE: b_i_k_6_i_j_0	// matmul/matmul-hw.mlir:14367:5
  assign c_prev_i_k_6_i_j_0 = C_reg_bank6_p0_rd_data_2447;	// matmul/matmul-hw.mlir:14213:31, :14369:5
  //PROBE: c_prev_i_k_6_i_j_0	// matmul/matmul-hw.mlir:14370:5
  assign tk_i_k_6_i_j_0 = _T_2775;	// matmul/matmul-hw.mlir:14372:5
  //PROBE: tk_i_k_6_i_j_0	// matmul/matmul-hw.mlir:14373:5
  wire [31:0] _T_2969 = mult_inst6_result + C_reg_bank6_p0_rd_data_2447;	// matmul/matmul-hw.mlir:14213:31, :14360:26, :14374:13
  assign c_i_k_6_i_j_0 = _T_2969;	// matmul/matmul-hw.mlir:14376:5
  //PROBE: c_i_k_6_i_j_0	// matmul/matmul-hw.mlir:14377:5
  assign _T_1355 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14378:13
  assign _T_1354 = _T_2819 ? _T_2969 : 32'bx;	// matmul/matmul-hw.mlir:9389:19, :14379:13
  assign _T_1353 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14380:13
  assign _T_1352 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14381:13
  mult mult_inst7 (	// matmul/matmul-hw.mlir:14382:26
    .a      (A_reg_bank7_p0_rd_data),	// matmul/matmul-hw.mlir:12222:31
    .b      (_T_2566),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst7_result)
  );
  assign _T_1351 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14383:13
  assign a_i_k_7_i_j_0 = A_reg_bank7_p0_rd_data;	// matmul/matmul-hw.mlir:12222:31, :14385:5
  //PROBE: a_i_k_7_i_j_0	// matmul/matmul-hw.mlir:14386:5
  assign b_i_k_7_i_j_0 = _T_2566;	// matmul/matmul-hw.mlir:14388:5
  //PROBE: b_i_k_7_i_j_0	// matmul/matmul-hw.mlir:14389:5
  assign c_prev_i_k_7_i_j_0 = C_reg_bank7_p0_rd_data_2446;	// matmul/matmul-hw.mlir:14214:31, :14391:5
  //PROBE: c_prev_i_k_7_i_j_0	// matmul/matmul-hw.mlir:14392:5
  assign tk_i_k_7_i_j_0 = _T_2786;	// matmul/matmul-hw.mlir:14394:5
  //PROBE: tk_i_k_7_i_j_0	// matmul/matmul-hw.mlir:14395:5
  wire [31:0] _T_2970 = mult_inst7_result + C_reg_bank7_p0_rd_data_2446;	// matmul/matmul-hw.mlir:14214:31, :14382:26, :14396:13
  assign c_i_k_7_i_j_0 = _T_2970;	// matmul/matmul-hw.mlir:14398:5
  //PROBE: c_i_k_7_i_j_0	// matmul/matmul-hw.mlir:14399:5
  assign _T_1350 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14400:13
  assign _T_1349 = _T_2830 ? _T_2970 : 32'bx;	// matmul/matmul-hw.mlir:9384:19, :14401:13
  assign _T_1348 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14402:13
  assign _T_1347 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14403:13
  mult mult_inst8 (	// matmul/matmul-hw.mlir:14404:26
    .a      (A_reg_bank8_p0_rd_data),	// matmul/matmul-hw.mlir:12223:31
    .b      (_T_2582),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst8_result)
  );
  assign _T_1346 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14405:13
  assign a_i_k_8_i_j_0 = A_reg_bank8_p0_rd_data;	// matmul/matmul-hw.mlir:12223:31, :14407:5
  //PROBE: a_i_k_8_i_j_0	// matmul/matmul-hw.mlir:14408:5
  assign b_i_k_8_i_j_0 = _T_2582;	// matmul/matmul-hw.mlir:14410:5
  //PROBE: b_i_k_8_i_j_0	// matmul/matmul-hw.mlir:14411:5
  assign c_prev_i_k_8_i_j_0 = C_reg_bank8_p0_rd_data_2445;	// matmul/matmul-hw.mlir:14215:31, :14413:5
  //PROBE: c_prev_i_k_8_i_j_0	// matmul/matmul-hw.mlir:14414:5
  assign tk_i_k_8_i_j_0 = _T_2797;	// matmul/matmul-hw.mlir:14416:5
  //PROBE: tk_i_k_8_i_j_0	// matmul/matmul-hw.mlir:14417:5
  wire [31:0] _T_2971 = mult_inst8_result + C_reg_bank8_p0_rd_data_2445;	// matmul/matmul-hw.mlir:14215:31, :14404:26, :14418:13
  assign c_i_k_8_i_j_0 = _T_2971;	// matmul/matmul-hw.mlir:14420:5
  //PROBE: c_i_k_8_i_j_0	// matmul/matmul-hw.mlir:14421:5
  assign _T_1345 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14422:13
  assign _T_1344 = _T_2841 ? _T_2971 : 32'bx;	// matmul/matmul-hw.mlir:9379:19, :14423:13
  assign _T_1343 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14424:13
  assign _T_1342 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14425:13
  mult mult_inst9 (	// matmul/matmul-hw.mlir:14426:26
    .a      (A_reg_bank9_p0_rd_data),	// matmul/matmul-hw.mlir:12224:31
    .b      (_T_2598),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst9_result)
  );
  assign _T_1341 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14427:13
  assign a_i_k_9_i_j_0 = A_reg_bank9_p0_rd_data;	// matmul/matmul-hw.mlir:12224:31, :14429:5
  //PROBE: a_i_k_9_i_j_0	// matmul/matmul-hw.mlir:14430:5
  assign b_i_k_9_i_j_0 = _T_2598;	// matmul/matmul-hw.mlir:14432:5
  //PROBE: b_i_k_9_i_j_0	// matmul/matmul-hw.mlir:14433:5
  assign c_prev_i_k_9_i_j_0 = C_reg_bank9_p0_rd_data_2444;	// matmul/matmul-hw.mlir:14216:31, :14435:5
  //PROBE: c_prev_i_k_9_i_j_0	// matmul/matmul-hw.mlir:14436:5
  assign tk_i_k_9_i_j_0 = _T_2808;	// matmul/matmul-hw.mlir:14438:5
  //PROBE: tk_i_k_9_i_j_0	// matmul/matmul-hw.mlir:14439:5
  wire [31:0] _T_2972 = mult_inst9_result + C_reg_bank9_p0_rd_data_2444;	// matmul/matmul-hw.mlir:14216:31, :14426:26, :14440:13
  assign c_i_k_9_i_j_0 = _T_2972;	// matmul/matmul-hw.mlir:14442:5
  //PROBE: c_i_k_9_i_j_0	// matmul/matmul-hw.mlir:14443:5
  assign _T_1340 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14444:13
  assign _T_1339 = _T_2852 ? _T_2972 : 32'bx;	// matmul/matmul-hw.mlir:9374:19, :14445:13
  assign _T_1338 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14446:13
  assign _T_1337 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14447:13
  mult mult_inst10 (	// matmul/matmul-hw.mlir:14448:27
    .a      (A_reg_bank10_p0_rd_data),	// matmul/matmul-hw.mlir:12225:32
    .b      (_T_2614),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst10_result)
  );
  assign _T_1336 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14449:13
  assign a_i_k_10_i_j_0 = A_reg_bank10_p0_rd_data;	// matmul/matmul-hw.mlir:12225:32, :14451:5
  //PROBE: a_i_k_10_i_j_0	// matmul/matmul-hw.mlir:14452:5
  assign b_i_k_10_i_j_0 = _T_2614;	// matmul/matmul-hw.mlir:14454:5
  //PROBE: b_i_k_10_i_j_0	// matmul/matmul-hw.mlir:14455:5
  assign c_prev_i_k_10_i_j_0 = C_reg_bank10_p0_rd_data_2443;	// matmul/matmul-hw.mlir:14217:32, :14457:5
  //PROBE: c_prev_i_k_10_i_j_0	// matmul/matmul-hw.mlir:14458:5
  assign tk_i_k_10_i_j_0 = _T_2819;	// matmul/matmul-hw.mlir:14460:5
  //PROBE: tk_i_k_10_i_j_0	// matmul/matmul-hw.mlir:14461:5
  wire [31:0] _T_2973 = mult_inst10_result + C_reg_bank10_p0_rd_data_2443;	// matmul/matmul-hw.mlir:14217:32, :14448:27, :14462:13
  assign c_i_k_10_i_j_0 = _T_2973;	// matmul/matmul-hw.mlir:14464:5
  //PROBE: c_i_k_10_i_j_0	// matmul/matmul-hw.mlir:14465:5
  assign _T_1335 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14466:13
  assign _T_1334 = _T_2863 ? _T_2973 : 32'bx;	// matmul/matmul-hw.mlir:9369:19, :14467:13
  assign _T_1333 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14468:13
  assign _T_1332 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14469:13
  mult mult_inst11 (	// matmul/matmul-hw.mlir:14470:27
    .a      (A_reg_bank11_p0_rd_data),	// matmul/matmul-hw.mlir:12226:32
    .b      (_T_2630),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst11_result)
  );
  assign _T_1331 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14471:13
  assign a_i_k_11_i_j_0 = A_reg_bank11_p0_rd_data;	// matmul/matmul-hw.mlir:12226:32, :14473:5
  //PROBE: a_i_k_11_i_j_0	// matmul/matmul-hw.mlir:14474:5
  assign b_i_k_11_i_j_0 = _T_2630;	// matmul/matmul-hw.mlir:14476:5
  //PROBE: b_i_k_11_i_j_0	// matmul/matmul-hw.mlir:14477:5
  assign c_prev_i_k_11_i_j_0 = C_reg_bank11_p0_rd_data_2442;	// matmul/matmul-hw.mlir:14218:32, :14479:5
  //PROBE: c_prev_i_k_11_i_j_0	// matmul/matmul-hw.mlir:14480:5
  assign tk_i_k_11_i_j_0 = _T_2830;	// matmul/matmul-hw.mlir:14482:5
  //PROBE: tk_i_k_11_i_j_0	// matmul/matmul-hw.mlir:14483:5
  wire [31:0] _T_2974 = mult_inst11_result + C_reg_bank11_p0_rd_data_2442;	// matmul/matmul-hw.mlir:14218:32, :14470:27, :14484:13
  assign c_i_k_11_i_j_0 = _T_2974;	// matmul/matmul-hw.mlir:14486:5
  //PROBE: c_i_k_11_i_j_0	// matmul/matmul-hw.mlir:14487:5
  assign _T_1330 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14488:13
  assign _T_1329 = _T_2874 ? _T_2974 : 32'bx;	// matmul/matmul-hw.mlir:9364:19, :14489:13
  assign _T_1328 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14490:13
  assign _T_1327 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14491:13
  mult mult_inst12 (	// matmul/matmul-hw.mlir:14492:27
    .a      (A_reg_bank12_p0_rd_data),	// matmul/matmul-hw.mlir:12227:32
    .b      (_T_2646),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst12_result)
  );
  assign _T_1326 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14493:13
  assign a_i_k_12_i_j_0 = A_reg_bank12_p0_rd_data;	// matmul/matmul-hw.mlir:12227:32, :14495:5
  //PROBE: a_i_k_12_i_j_0	// matmul/matmul-hw.mlir:14496:5
  assign b_i_k_12_i_j_0 = _T_2646;	// matmul/matmul-hw.mlir:14498:5
  //PROBE: b_i_k_12_i_j_0	// matmul/matmul-hw.mlir:14499:5
  assign c_prev_i_k_12_i_j_0 = C_reg_bank12_p0_rd_data_2441;	// matmul/matmul-hw.mlir:14219:32, :14501:5
  //PROBE: c_prev_i_k_12_i_j_0	// matmul/matmul-hw.mlir:14502:5
  assign tk_i_k_12_i_j_0 = _T_2841;	// matmul/matmul-hw.mlir:14504:5
  //PROBE: tk_i_k_12_i_j_0	// matmul/matmul-hw.mlir:14505:5
  wire [31:0] _T_2975 = mult_inst12_result + C_reg_bank12_p0_rd_data_2441;	// matmul/matmul-hw.mlir:14219:32, :14492:27, :14506:13
  assign c_i_k_12_i_j_0 = _T_2975;	// matmul/matmul-hw.mlir:14508:5
  //PROBE: c_i_k_12_i_j_0	// matmul/matmul-hw.mlir:14509:5
  assign _T_1325 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14510:13
  assign _T_1324 = _T_2885 ? _T_2975 : 32'bx;	// matmul/matmul-hw.mlir:9359:19, :14511:13
  assign _T_1323 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14512:13
  assign _T_1322 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14513:13
  mult mult_inst13 (	// matmul/matmul-hw.mlir:14514:27
    .a      (A_reg_bank13_p0_rd_data),	// matmul/matmul-hw.mlir:12228:32
    .b      (_T_2662),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst13_result)
  );
  assign _T_1321 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14515:13
  assign a_i_k_13_i_j_0 = A_reg_bank13_p0_rd_data;	// matmul/matmul-hw.mlir:12228:32, :14517:5
  //PROBE: a_i_k_13_i_j_0	// matmul/matmul-hw.mlir:14518:5
  assign b_i_k_13_i_j_0 = _T_2662;	// matmul/matmul-hw.mlir:14520:5
  //PROBE: b_i_k_13_i_j_0	// matmul/matmul-hw.mlir:14521:5
  assign c_prev_i_k_13_i_j_0 = C_reg_bank13_p0_rd_data_2440;	// matmul/matmul-hw.mlir:14220:32, :14523:5
  //PROBE: c_prev_i_k_13_i_j_0	// matmul/matmul-hw.mlir:14524:5
  assign tk_i_k_13_i_j_0 = _T_2852;	// matmul/matmul-hw.mlir:14526:5
  //PROBE: tk_i_k_13_i_j_0	// matmul/matmul-hw.mlir:14527:5
  wire [31:0] _T_2976 = mult_inst13_result + C_reg_bank13_p0_rd_data_2440;	// matmul/matmul-hw.mlir:14220:32, :14514:27, :14528:13
  assign c_i_k_13_i_j_0 = _T_2976;	// matmul/matmul-hw.mlir:14530:5
  //PROBE: c_i_k_13_i_j_0	// matmul/matmul-hw.mlir:14531:5
  assign _T_1320 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14532:13
  assign _T_1319 = _T_2892 ? _T_2976 : 32'bx;	// matmul/matmul-hw.mlir:9354:19, :14533:13
  assign _T_1318 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14534:13
  assign _T_1317 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14535:13
  mult mult_inst14 (	// matmul/matmul-hw.mlir:14536:27
    .a      (A_reg_bank14_p0_rd_data),	// matmul/matmul-hw.mlir:12229:32
    .b      (_T_2678),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst14_result)
  );
  assign _T_1316 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14537:13
  assign a_i_k_14_i_j_0 = A_reg_bank14_p0_rd_data;	// matmul/matmul-hw.mlir:12229:32, :14539:5
  //PROBE: a_i_k_14_i_j_0	// matmul/matmul-hw.mlir:14540:5
  assign b_i_k_14_i_j_0 = _T_2678;	// matmul/matmul-hw.mlir:14542:5
  //PROBE: b_i_k_14_i_j_0	// matmul/matmul-hw.mlir:14543:5
  assign c_prev_i_k_14_i_j_0 = C_reg_bank14_p0_rd_data_2439;	// matmul/matmul-hw.mlir:14221:32, :14545:5
  //PROBE: c_prev_i_k_14_i_j_0	// matmul/matmul-hw.mlir:14546:5
  assign tk_i_k_14_i_j_0 = _T_2863;	// matmul/matmul-hw.mlir:14548:5
  //PROBE: tk_i_k_14_i_j_0	// matmul/matmul-hw.mlir:14549:5
  wire [31:0] _T_2977 = mult_inst14_result + C_reg_bank14_p0_rd_data_2439;	// matmul/matmul-hw.mlir:14221:32, :14536:27, :14550:13
  assign c_i_k_14_i_j_0 = _T_2977;	// matmul/matmul-hw.mlir:14552:5
  //PROBE: c_i_k_14_i_j_0	// matmul/matmul-hw.mlir:14553:5
  assign _T_1315 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14554:13
  assign _T_1314 = _T_2897 ? _T_2977 : 32'bx;	// matmul/matmul-hw.mlir:9349:19, :14555:13
  assign _T_1313 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14556:13
  assign _T_1312 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14557:13
  mult mult_inst15 (	// matmul/matmul-hw.mlir:14558:27
    .a      (A_reg_bank15_p0_rd_data),	// matmul/matmul-hw.mlir:12230:32
    .b      (_T_2694),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst15_result)
  );
  assign _T_1311 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14559:13
  assign a_i_k_15_i_j_0 = A_reg_bank15_p0_rd_data;	// matmul/matmul-hw.mlir:12230:32, :14561:5
  //PROBE: a_i_k_15_i_j_0	// matmul/matmul-hw.mlir:14562:5
  assign b_i_k_15_i_j_0 = _T_2694;	// matmul/matmul-hw.mlir:14564:5
  //PROBE: b_i_k_15_i_j_0	// matmul/matmul-hw.mlir:14565:5
  assign c_prev_i_k_15_i_j_0 = C_reg_bank15_p0_rd_data_2438;	// matmul/matmul-hw.mlir:14222:32, :14567:5
  //PROBE: c_prev_i_k_15_i_j_0	// matmul/matmul-hw.mlir:14568:5
  assign tk_i_k_15_i_j_0 = _T_2874;	// matmul/matmul-hw.mlir:14570:5
  //PROBE: tk_i_k_15_i_j_0	// matmul/matmul-hw.mlir:14571:5
  wire [31:0] _T_2978 = mult_inst15_result + C_reg_bank15_p0_rd_data_2438;	// matmul/matmul-hw.mlir:14222:32, :14558:27, :14572:13
  assign c_i_k_15_i_j_0 = _T_2978;	// matmul/matmul-hw.mlir:14574:5
  //PROBE: c_i_k_15_i_j_0	// matmul/matmul-hw.mlir:14575:5
  assign _T_1310 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14576:13
  assign _T_1309 = _T_2902 ? _T_2978 : 32'bx;	// matmul/matmul-hw.mlir:9344:19, :14577:13
  assign _T_1308 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14578:13
  wire [3:0][3:0] _T_2979 = i_delayed;	// matmul/matmul-hw.mlir:14580:13
  wire [3:0][3:0] _T_2980 = {_T_2979[2'h0+:3], {{i_k_next_2886}}};	// matmul/matmul-hw.mlir:13184:12, :14581:19, :14582:13, :14583:13, :14584:13
  wire [3:0][3:0] _T_2981 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:14585:19, :14586:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14587:5
    if (rst)	// matmul/matmul-hw.mlir:14587:5
      i_delayed <= _T_2981;	// matmul/matmul-hw.mlir:14590:7
    else	// matmul/matmul-hw.mlir:14587:5
      i_delayed <= _T_2980;	// matmul/matmul-hw.mlir:14588:7
  end // always @(posedge)
  assign _T_1307 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14594:13
  assign _T_1306 = _T_2907 ? i_delayed[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:9341:18, :14580:13, :14592:20, :14593:13, :14595:13
  assign _T_1305 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14596:13
  assign _T_1304 = _T_2907 ? C_reg_bank16_p0_rd_data_2437 : 32'bx;	// matmul/matmul-hw.mlir:9339:19, :14223:32, :14597:13
  localparam [3:0] _T_2982 = 4'h0;	// matmul/matmul-hw.mlir:14600:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14601:5
    if (rst)	// matmul/matmul-hw.mlir:14601:5
      i_j_next <= _T_2982;	// matmul/matmul-hw.mlir:14604:7
    else	// matmul/matmul-hw.mlir:14601:5
      i_j_next <= _T_2718;	// matmul/matmul-hw.mlir:14602:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_2983 (	// matmul/matmul-hw.mlir:14674:36
    .p0_rd_en   (_T_1299),	// matmul/matmul-hw.mlir:14696:13
    .p1_wr_en   (_T_1303),	// matmul/matmul-hw.mlir:14691:13
    .p1_wr_data (_T_1302),	// matmul/matmul-hw.mlir:14692:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2436)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_2984 (	// matmul/matmul-hw.mlir:14675:36
    .p0_rd_en   (_T_1294),	// matmul/matmul-hw.mlir:14726:13
    .p1_wr_en   (_T_1298),	// matmul/matmul-hw.mlir:14713:13
    .p1_wr_data (_T_1297),	// matmul/matmul-hw.mlir:14714:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2435)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_2985 (	// matmul/matmul-hw.mlir:14676:36
    .p0_rd_en   (_T_1289),	// matmul/matmul-hw.mlir:14756:13
    .p1_wr_en   (_T_1293),	// matmul/matmul-hw.mlir:14743:13
    .p1_wr_data (_T_1292),	// matmul/matmul-hw.mlir:14744:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2434)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_2986 (	// matmul/matmul-hw.mlir:14677:36
    .p0_rd_en   (_T_1284),	// matmul/matmul-hw.mlir:14786:13
    .p1_wr_en   (_T_1288),	// matmul/matmul-hw.mlir:14773:13
    .p1_wr_data (_T_1287),	// matmul/matmul-hw.mlir:14774:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2433)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_2987 (	// matmul/matmul-hw.mlir:14678:36
    .p0_rd_en   (_T_1279),	// matmul/matmul-hw.mlir:14816:13
    .p1_wr_en   (_T_1283),	// matmul/matmul-hw.mlir:14803:13
    .p1_wr_data (_T_1282),	// matmul/matmul-hw.mlir:14804:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2432)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_2988 (	// matmul/matmul-hw.mlir:14679:36
    .p0_rd_en   (_T_1274),	// matmul/matmul-hw.mlir:14846:13
    .p1_wr_en   (_T_1278),	// matmul/matmul-hw.mlir:14833:13
    .p1_wr_data (_T_1277),	// matmul/matmul-hw.mlir:14834:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2431)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_2989 (	// matmul/matmul-hw.mlir:14680:36
    .p0_rd_en   (_T_1269),	// matmul/matmul-hw.mlir:14876:13
    .p1_wr_en   (_T_1273),	// matmul/matmul-hw.mlir:14863:13
    .p1_wr_data (_T_1272),	// matmul/matmul-hw.mlir:14864:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2430)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_2990 (	// matmul/matmul-hw.mlir:14681:36
    .p0_rd_en   (_T_1264),	// matmul/matmul-hw.mlir:14906:13
    .p1_wr_en   (_T_1268),	// matmul/matmul-hw.mlir:14893:13
    .p1_wr_data (_T_1267),	// matmul/matmul-hw.mlir:14894:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2429)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_2991 (	// matmul/matmul-hw.mlir:14682:36
    .p0_rd_en   (_T_1259),	// matmul/matmul-hw.mlir:14936:13
    .p1_wr_en   (_T_1263),	// matmul/matmul-hw.mlir:14923:13
    .p1_wr_data (_T_1262),	// matmul/matmul-hw.mlir:14924:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2428)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_2992 (	// matmul/matmul-hw.mlir:14683:36
    .p0_rd_en   (_T_1254),	// matmul/matmul-hw.mlir:14966:13
    .p1_wr_en   (_T_1258),	// matmul/matmul-hw.mlir:14953:13
    .p1_wr_data (_T_1257),	// matmul/matmul-hw.mlir:14954:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2427)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_2993 (	// matmul/matmul-hw.mlir:14684:37
    .p0_rd_en   (_T_1249),	// matmul/matmul-hw.mlir:14996:13
    .p1_wr_en   (_T_1253),	// matmul/matmul-hw.mlir:14983:13
    .p1_wr_data (_T_1252),	// matmul/matmul-hw.mlir:14984:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2426)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_2994 (	// matmul/matmul-hw.mlir:14685:37
    .p0_rd_en   (_T_1244),	// matmul/matmul-hw.mlir:15026:13
    .p1_wr_en   (_T_1248),	// matmul/matmul-hw.mlir:15013:13
    .p1_wr_data (_T_1247),	// matmul/matmul-hw.mlir:15014:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2425)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_2995 (	// matmul/matmul-hw.mlir:14686:37
    .p0_rd_en   (_T_1239),	// matmul/matmul-hw.mlir:15056:13
    .p1_wr_en   (_T_1243),	// matmul/matmul-hw.mlir:15043:13
    .p1_wr_data (_T_1242),	// matmul/matmul-hw.mlir:15044:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2424)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_2996 (	// matmul/matmul-hw.mlir:14687:37
    .p0_rd_en   (_T_1234),	// matmul/matmul-hw.mlir:15086:13
    .p1_wr_en   (_T_1238),	// matmul/matmul-hw.mlir:15073:13
    .p1_wr_data (_T_1237),	// matmul/matmul-hw.mlir:15074:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2423)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_2997 (	// matmul/matmul-hw.mlir:14688:37
    .p0_rd_en   (_T_1229),	// matmul/matmul-hw.mlir:15116:13
    .p1_wr_en   (_T_1233),	// matmul/matmul-hw.mlir:15103:13
    .p1_wr_data (_T_1232),	// matmul/matmul-hw.mlir:15104:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2422)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_2998 (	// matmul/matmul-hw.mlir:14689:37
    .p0_rd_en   (_T_1224),	// matmul/matmul-hw.mlir:15146:13
    .p1_wr_en   (_T_1228),	// matmul/matmul-hw.mlir:15133:13
    .p1_wr_data (_T_1227),	// matmul/matmul-hw.mlir:15134:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2421)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_2999 (	// matmul/matmul-hw.mlir:14690:37
    .p0_rd_en   (_T_1221),	// matmul/matmul-hw.mlir:15173:13
    .p1_wr_en   (_T_1223),	// matmul/matmul-hw.mlir:15163:13
    .p1_wr_data (_T_1222),	// matmul/matmul-hw.mlir:15164:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2420)
  );
  assign _T_1303 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14691:13
  assign _T_1302 = _T_2753 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :9337:19, :14692:13
  assign _T_1301 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14693:13
  assign _T_1300 = _T_2742 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14694:13
  mult mult_inst16 (	// matmul/matmul-hw.mlir:14695:27
    .a      (A_reg_bank16_p0_rd_data),	// matmul/matmul-hw.mlir:12231:32
    .b      (_T_2455),
    .t      (_T_2742),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst16_result)
  );
  assign _T_1299 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14696:13
  assign a_i_k_0_i_j_1 = A_reg_bank16_p0_rd_data;	// matmul/matmul-hw.mlir:12231:32, :14698:5
  //PROBE: a_i_k_0_i_j_1	// matmul/matmul-hw.mlir:14699:5
  assign b_i_k_0_i_j_1 = _T_2455;	// matmul/matmul-hw.mlir:14701:5
  //PROBE: b_i_k_0_i_j_1	// matmul/matmul-hw.mlir:14702:5
  assign c_prev_i_k_0_i_j_1 = C_reg_bank0_p0_rd_data_2436;	// matmul/matmul-hw.mlir:14674:36, :14704:5
  //PROBE: c_prev_i_k_0_i_j_1	// matmul/matmul-hw.mlir:14705:5
  assign tk_i_k_0_i_j_1 = _T_2189;	// matmul/matmul-hw.mlir:12484:12, :14707:5
  //PROBE: tk_i_k_0_i_j_1	// matmul/matmul-hw.mlir:14708:5
  wire [31:0] _T_3000 = mult_inst16_result + C_reg_bank0_p0_rd_data_2436;	// matmul/matmul-hw.mlir:14674:36, :14695:27, :14709:13
  assign c_i_k_0_i_j_1 = _T_3000;	// matmul/matmul-hw.mlir:14711:5
  //PROBE: c_i_k_0_i_j_1	// matmul/matmul-hw.mlir:14712:5
  assign _T_1298 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14713:13
  assign _T_1297 = _T_2764 ? _T_3000 : 32'bx;	// matmul/matmul-hw.mlir:9332:19, :14714:13
  localparam [3:0] _T_3002 = 4'h0;	// matmul/matmul-hw.mlir:14717:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14718:5
    if (rst)	// matmul/matmul-hw.mlir:14718:5
      i_k_next_3001 <= _T_3002;	// matmul/matmul-hw.mlir:14721:7
    else	// matmul/matmul-hw.mlir:14718:5
      i_k_next_3001 <= i_j_next;	// matmul/matmul-hw.mlir:14599:13, :14719:7
  end // always @(posedge)
  assign _T_1296 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14723:13
  assign _T_1295 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14724:13
  mult mult_inst17 (	// matmul/matmul-hw.mlir:14725:27
    .a      (A_reg_bank17_p0_rd_data),	// matmul/matmul-hw.mlir:12232:32
    .b      (_T_2471),
    .t      (_T_2753),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst17_result)
  );
  assign _T_1294 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14726:13
  assign a_i_k_1_i_j_1 = A_reg_bank17_p0_rd_data;	// matmul/matmul-hw.mlir:12232:32, :14728:5
  //PROBE: a_i_k_1_i_j_1	// matmul/matmul-hw.mlir:14729:5
  assign b_i_k_1_i_j_1 = _T_2471;	// matmul/matmul-hw.mlir:14731:5
  //PROBE: b_i_k_1_i_j_1	// matmul/matmul-hw.mlir:14732:5
  assign c_prev_i_k_1_i_j_1 = C_reg_bank1_p0_rd_data_2435;	// matmul/matmul-hw.mlir:14675:36, :14734:5
  //PROBE: c_prev_i_k_1_i_j_1	// matmul/matmul-hw.mlir:14735:5
  assign tk_i_k_1_i_j_1 = _T_2731;	// matmul/matmul-hw.mlir:14737:5
  //PROBE: tk_i_k_1_i_j_1	// matmul/matmul-hw.mlir:14738:5
  wire [31:0] _T_3003 = mult_inst17_result + C_reg_bank1_p0_rd_data_2435;	// matmul/matmul-hw.mlir:14675:36, :14725:27, :14739:13
  assign c_i_k_1_i_j_1 = _T_3003;	// matmul/matmul-hw.mlir:14741:5
  //PROBE: c_i_k_1_i_j_1	// matmul/matmul-hw.mlir:14742:5
  assign _T_1293 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14743:13
  assign _T_1292 = _T_2775 ? _T_3003 : 32'bx;	// matmul/matmul-hw.mlir:9327:19, :14744:13
  localparam [3:0] _T_3005 = 4'h0;	// matmul/matmul-hw.mlir:14747:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14748:5
    if (rst)	// matmul/matmul-hw.mlir:14748:5
      i_k_next_3004 <= _T_3005;	// matmul/matmul-hw.mlir:14751:7
    else	// matmul/matmul-hw.mlir:14748:5
      i_k_next_3004 <= i_k_next_3001;	// matmul/matmul-hw.mlir:14716:13, :14749:7
  end // always @(posedge)
  assign _T_1291 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14753:13
  assign _T_1290 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14754:13
  mult mult_inst18 (	// matmul/matmul-hw.mlir:14755:27
    .a      (A_reg_bank18_p0_rd_data),	// matmul/matmul-hw.mlir:12233:32
    .b      (_T_2487),
    .t      (_T_2764),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst18_result)
  );
  assign _T_1289 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14756:13
  assign a_i_k_2_i_j_1 = A_reg_bank18_p0_rd_data;	// matmul/matmul-hw.mlir:12233:32, :14758:5
  //PROBE: a_i_k_2_i_j_1	// matmul/matmul-hw.mlir:14759:5
  assign b_i_k_2_i_j_1 = _T_2487;	// matmul/matmul-hw.mlir:14761:5
  //PROBE: b_i_k_2_i_j_1	// matmul/matmul-hw.mlir:14762:5
  assign c_prev_i_k_2_i_j_1 = C_reg_bank2_p0_rd_data_2434;	// matmul/matmul-hw.mlir:14676:36, :14764:5
  //PROBE: c_prev_i_k_2_i_j_1	// matmul/matmul-hw.mlir:14765:5
  assign tk_i_k_2_i_j_1 = _T_2742;	// matmul/matmul-hw.mlir:14767:5
  //PROBE: tk_i_k_2_i_j_1	// matmul/matmul-hw.mlir:14768:5
  wire [31:0] _T_3006 = mult_inst18_result + C_reg_bank2_p0_rd_data_2434;	// matmul/matmul-hw.mlir:14676:36, :14755:27, :14769:13
  assign c_i_k_2_i_j_1 = _T_3006;	// matmul/matmul-hw.mlir:14771:5
  //PROBE: c_i_k_2_i_j_1	// matmul/matmul-hw.mlir:14772:5
  assign _T_1288 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14773:13
  assign _T_1287 = _T_2786 ? _T_3006 : 32'bx;	// matmul/matmul-hw.mlir:9322:19, :14774:13
  localparam [3:0] _T_3008 = 4'h0;	// matmul/matmul-hw.mlir:14777:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14778:5
    if (rst)	// matmul/matmul-hw.mlir:14778:5
      i_k_next_3007 <= _T_3008;	// matmul/matmul-hw.mlir:14781:7
    else	// matmul/matmul-hw.mlir:14778:5
      i_k_next_3007 <= i_k_next_3004;	// matmul/matmul-hw.mlir:14746:13, :14779:7
  end // always @(posedge)
  assign _T_1286 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14783:13
  assign _T_1285 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14784:13
  mult mult_inst19 (	// matmul/matmul-hw.mlir:14785:27
    .a      (A_reg_bank19_p0_rd_data),	// matmul/matmul-hw.mlir:12234:32
    .b      (_T_2503),
    .t      (_T_2775),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst19_result)
  );
  assign _T_1284 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14786:13
  assign a_i_k_3_i_j_1 = A_reg_bank19_p0_rd_data;	// matmul/matmul-hw.mlir:12234:32, :14788:5
  //PROBE: a_i_k_3_i_j_1	// matmul/matmul-hw.mlir:14789:5
  assign b_i_k_3_i_j_1 = _T_2503;	// matmul/matmul-hw.mlir:14791:5
  //PROBE: b_i_k_3_i_j_1	// matmul/matmul-hw.mlir:14792:5
  assign c_prev_i_k_3_i_j_1 = C_reg_bank3_p0_rd_data_2433;	// matmul/matmul-hw.mlir:14677:36, :14794:5
  //PROBE: c_prev_i_k_3_i_j_1	// matmul/matmul-hw.mlir:14795:5
  assign tk_i_k_3_i_j_1 = _T_2753;	// matmul/matmul-hw.mlir:14797:5
  //PROBE: tk_i_k_3_i_j_1	// matmul/matmul-hw.mlir:14798:5
  wire [31:0] _T_3009 = mult_inst19_result + C_reg_bank3_p0_rd_data_2433;	// matmul/matmul-hw.mlir:14677:36, :14785:27, :14799:13
  assign c_i_k_3_i_j_1 = _T_3009;	// matmul/matmul-hw.mlir:14801:5
  //PROBE: c_i_k_3_i_j_1	// matmul/matmul-hw.mlir:14802:5
  assign _T_1283 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14803:13
  assign _T_1282 = _T_2797 ? _T_3009 : 32'bx;	// matmul/matmul-hw.mlir:9317:19, :14804:13
  localparam [3:0] _T_3011 = 4'h0;	// matmul/matmul-hw.mlir:14807:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14808:5
    if (rst)	// matmul/matmul-hw.mlir:14808:5
      i_k_next_3010 <= _T_3011;	// matmul/matmul-hw.mlir:14811:7
    else	// matmul/matmul-hw.mlir:14808:5
      i_k_next_3010 <= i_k_next_3007;	// matmul/matmul-hw.mlir:14776:13, :14809:7
  end // always @(posedge)
  assign _T_1281 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14813:13
  assign _T_1280 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14814:13
  mult mult_inst20 (	// matmul/matmul-hw.mlir:14815:27
    .a      (A_reg_bank20_p0_rd_data),	// matmul/matmul-hw.mlir:12235:32
    .b      (_T_2519),
    .t      (_T_2786),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst20_result)
  );
  assign _T_1279 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14816:13
  assign a_i_k_4_i_j_1 = A_reg_bank20_p0_rd_data;	// matmul/matmul-hw.mlir:12235:32, :14818:5
  //PROBE: a_i_k_4_i_j_1	// matmul/matmul-hw.mlir:14819:5
  assign b_i_k_4_i_j_1 = _T_2519;	// matmul/matmul-hw.mlir:14821:5
  //PROBE: b_i_k_4_i_j_1	// matmul/matmul-hw.mlir:14822:5
  assign c_prev_i_k_4_i_j_1 = C_reg_bank4_p0_rd_data_2432;	// matmul/matmul-hw.mlir:14678:36, :14824:5
  //PROBE: c_prev_i_k_4_i_j_1	// matmul/matmul-hw.mlir:14825:5
  assign tk_i_k_4_i_j_1 = _T_2764;	// matmul/matmul-hw.mlir:14827:5
  //PROBE: tk_i_k_4_i_j_1	// matmul/matmul-hw.mlir:14828:5
  wire [31:0] _T_3012 = mult_inst20_result + C_reg_bank4_p0_rd_data_2432;	// matmul/matmul-hw.mlir:14678:36, :14815:27, :14829:13
  assign c_i_k_4_i_j_1 = _T_3012;	// matmul/matmul-hw.mlir:14831:5
  //PROBE: c_i_k_4_i_j_1	// matmul/matmul-hw.mlir:14832:5
  assign _T_1278 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14833:13
  assign _T_1277 = _T_2808 ? _T_3012 : 32'bx;	// matmul/matmul-hw.mlir:9312:19, :14834:13
  localparam [3:0] _T_3014 = 4'h0;	// matmul/matmul-hw.mlir:14837:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14838:5
    if (rst)	// matmul/matmul-hw.mlir:14838:5
      i_k_next_3013 <= _T_3014;	// matmul/matmul-hw.mlir:14841:7
    else	// matmul/matmul-hw.mlir:14838:5
      i_k_next_3013 <= i_k_next_3010;	// matmul/matmul-hw.mlir:14806:13, :14839:7
  end // always @(posedge)
  assign _T_1276 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14843:13
  assign _T_1275 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14844:13
  mult mult_inst21 (	// matmul/matmul-hw.mlir:14845:27
    .a      (A_reg_bank21_p0_rd_data),	// matmul/matmul-hw.mlir:12236:32
    .b      (_T_2535),
    .t      (_T_2797),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst21_result)
  );
  assign _T_1274 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14846:13
  assign a_i_k_5_i_j_1 = A_reg_bank21_p0_rd_data;	// matmul/matmul-hw.mlir:12236:32, :14848:5
  //PROBE: a_i_k_5_i_j_1	// matmul/matmul-hw.mlir:14849:5
  assign b_i_k_5_i_j_1 = _T_2535;	// matmul/matmul-hw.mlir:14851:5
  //PROBE: b_i_k_5_i_j_1	// matmul/matmul-hw.mlir:14852:5
  assign c_prev_i_k_5_i_j_1 = C_reg_bank5_p0_rd_data_2431;	// matmul/matmul-hw.mlir:14679:36, :14854:5
  //PROBE: c_prev_i_k_5_i_j_1	// matmul/matmul-hw.mlir:14855:5
  assign tk_i_k_5_i_j_1 = _T_2775;	// matmul/matmul-hw.mlir:14857:5
  //PROBE: tk_i_k_5_i_j_1	// matmul/matmul-hw.mlir:14858:5
  wire [31:0] _T_3015 = mult_inst21_result + C_reg_bank5_p0_rd_data_2431;	// matmul/matmul-hw.mlir:14679:36, :14845:27, :14859:13
  assign c_i_k_5_i_j_1 = _T_3015;	// matmul/matmul-hw.mlir:14861:5
  //PROBE: c_i_k_5_i_j_1	// matmul/matmul-hw.mlir:14862:5
  assign _T_1273 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14863:13
  assign _T_1272 = _T_2819 ? _T_3015 : 32'bx;	// matmul/matmul-hw.mlir:9307:19, :14864:13
  localparam [3:0] _T_3017 = 4'h0;	// matmul/matmul-hw.mlir:14867:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14868:5
    if (rst)	// matmul/matmul-hw.mlir:14868:5
      i_k_next_3016 <= _T_3017;	// matmul/matmul-hw.mlir:14871:7
    else	// matmul/matmul-hw.mlir:14868:5
      i_k_next_3016 <= i_k_next_3013;	// matmul/matmul-hw.mlir:14836:13, :14869:7
  end // always @(posedge)
  assign _T_1271 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14873:13
  assign _T_1270 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14874:13
  mult mult_inst22 (	// matmul/matmul-hw.mlir:14875:27
    .a      (A_reg_bank22_p0_rd_data),	// matmul/matmul-hw.mlir:12237:32
    .b      (_T_2551),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst22_result)
  );
  assign _T_1269 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14876:13
  assign a_i_k_6_i_j_1 = A_reg_bank22_p0_rd_data;	// matmul/matmul-hw.mlir:12237:32, :14878:5
  //PROBE: a_i_k_6_i_j_1	// matmul/matmul-hw.mlir:14879:5
  assign b_i_k_6_i_j_1 = _T_2551;	// matmul/matmul-hw.mlir:14881:5
  //PROBE: b_i_k_6_i_j_1	// matmul/matmul-hw.mlir:14882:5
  assign c_prev_i_k_6_i_j_1 = C_reg_bank6_p0_rd_data_2430;	// matmul/matmul-hw.mlir:14680:36, :14884:5
  //PROBE: c_prev_i_k_6_i_j_1	// matmul/matmul-hw.mlir:14885:5
  assign tk_i_k_6_i_j_1 = _T_2786;	// matmul/matmul-hw.mlir:14887:5
  //PROBE: tk_i_k_6_i_j_1	// matmul/matmul-hw.mlir:14888:5
  wire [31:0] _T_3018 = mult_inst22_result + C_reg_bank6_p0_rd_data_2430;	// matmul/matmul-hw.mlir:14680:36, :14875:27, :14889:13
  assign c_i_k_6_i_j_1 = _T_3018;	// matmul/matmul-hw.mlir:14891:5
  //PROBE: c_i_k_6_i_j_1	// matmul/matmul-hw.mlir:14892:5
  assign _T_1268 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14893:13
  assign _T_1267 = _T_2830 ? _T_3018 : 32'bx;	// matmul/matmul-hw.mlir:9302:19, :14894:13
  localparam [3:0] _T_3020 = 4'h0;	// matmul/matmul-hw.mlir:14897:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14898:5
    if (rst)	// matmul/matmul-hw.mlir:14898:5
      i_k_next_3019 <= _T_3020;	// matmul/matmul-hw.mlir:14901:7
    else	// matmul/matmul-hw.mlir:14898:5
      i_k_next_3019 <= i_k_next_3016;	// matmul/matmul-hw.mlir:14866:13, :14899:7
  end // always @(posedge)
  assign _T_1266 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14903:13
  assign _T_1265 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14904:13
  mult mult_inst23 (	// matmul/matmul-hw.mlir:14905:27
    .a      (A_reg_bank23_p0_rd_data),	// matmul/matmul-hw.mlir:12238:32
    .b      (_T_2567),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst23_result)
  );
  assign _T_1264 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14906:13
  assign a_i_k_7_i_j_1 = A_reg_bank23_p0_rd_data;	// matmul/matmul-hw.mlir:12238:32, :14908:5
  //PROBE: a_i_k_7_i_j_1	// matmul/matmul-hw.mlir:14909:5
  assign b_i_k_7_i_j_1 = _T_2567;	// matmul/matmul-hw.mlir:14911:5
  //PROBE: b_i_k_7_i_j_1	// matmul/matmul-hw.mlir:14912:5
  assign c_prev_i_k_7_i_j_1 = C_reg_bank7_p0_rd_data_2429;	// matmul/matmul-hw.mlir:14681:36, :14914:5
  //PROBE: c_prev_i_k_7_i_j_1	// matmul/matmul-hw.mlir:14915:5
  assign tk_i_k_7_i_j_1 = _T_2797;	// matmul/matmul-hw.mlir:14917:5
  //PROBE: tk_i_k_7_i_j_1	// matmul/matmul-hw.mlir:14918:5
  wire [31:0] _T_3021 = mult_inst23_result + C_reg_bank7_p0_rd_data_2429;	// matmul/matmul-hw.mlir:14681:36, :14905:27, :14919:13
  assign c_i_k_7_i_j_1 = _T_3021;	// matmul/matmul-hw.mlir:14921:5
  //PROBE: c_i_k_7_i_j_1	// matmul/matmul-hw.mlir:14922:5
  assign _T_1263 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14923:13
  assign _T_1262 = _T_2841 ? _T_3021 : 32'bx;	// matmul/matmul-hw.mlir:9297:19, :14924:13
  localparam [3:0] _T_3023 = 4'h0;	// matmul/matmul-hw.mlir:14927:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14928:5
    if (rst)	// matmul/matmul-hw.mlir:14928:5
      i_k_next_3022 <= _T_3023;	// matmul/matmul-hw.mlir:14931:7
    else	// matmul/matmul-hw.mlir:14928:5
      i_k_next_3022 <= i_k_next_3019;	// matmul/matmul-hw.mlir:14896:13, :14929:7
  end // always @(posedge)
  assign _T_1261 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14933:13
  assign _T_1260 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14934:13
  mult mult_inst24 (	// matmul/matmul-hw.mlir:14935:27
    .a      (A_reg_bank24_p0_rd_data),	// matmul/matmul-hw.mlir:12239:32
    .b      (_T_2583),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst24_result)
  );
  assign _T_1259 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14936:13
  assign a_i_k_8_i_j_1 = A_reg_bank24_p0_rd_data;	// matmul/matmul-hw.mlir:12239:32, :14938:5
  //PROBE: a_i_k_8_i_j_1	// matmul/matmul-hw.mlir:14939:5
  assign b_i_k_8_i_j_1 = _T_2583;	// matmul/matmul-hw.mlir:14941:5
  //PROBE: b_i_k_8_i_j_1	// matmul/matmul-hw.mlir:14942:5
  assign c_prev_i_k_8_i_j_1 = C_reg_bank8_p0_rd_data_2428;	// matmul/matmul-hw.mlir:14682:36, :14944:5
  //PROBE: c_prev_i_k_8_i_j_1	// matmul/matmul-hw.mlir:14945:5
  assign tk_i_k_8_i_j_1 = _T_2808;	// matmul/matmul-hw.mlir:14947:5
  //PROBE: tk_i_k_8_i_j_1	// matmul/matmul-hw.mlir:14948:5
  wire [31:0] _T_3024 = mult_inst24_result + C_reg_bank8_p0_rd_data_2428;	// matmul/matmul-hw.mlir:14682:36, :14935:27, :14949:13
  assign c_i_k_8_i_j_1 = _T_3024;	// matmul/matmul-hw.mlir:14951:5
  //PROBE: c_i_k_8_i_j_1	// matmul/matmul-hw.mlir:14952:5
  assign _T_1258 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14953:13
  assign _T_1257 = _T_2852 ? _T_3024 : 32'bx;	// matmul/matmul-hw.mlir:9292:19, :14954:13
  localparam [3:0] _T_3026 = 4'h0;	// matmul/matmul-hw.mlir:14957:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14958:5
    if (rst)	// matmul/matmul-hw.mlir:14958:5
      i_k_next_3025 <= _T_3026;	// matmul/matmul-hw.mlir:14961:7
    else	// matmul/matmul-hw.mlir:14958:5
      i_k_next_3025 <= i_k_next_3022;	// matmul/matmul-hw.mlir:14926:13, :14959:7
  end // always @(posedge)
  assign _T_1256 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14963:13
  assign _T_1255 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14964:13
  mult mult_inst25 (	// matmul/matmul-hw.mlir:14965:27
    .a      (A_reg_bank25_p0_rd_data),	// matmul/matmul-hw.mlir:12240:32
    .b      (_T_2599),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst25_result)
  );
  assign _T_1254 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14966:13
  assign a_i_k_9_i_j_1 = A_reg_bank25_p0_rd_data;	// matmul/matmul-hw.mlir:12240:32, :14968:5
  //PROBE: a_i_k_9_i_j_1	// matmul/matmul-hw.mlir:14969:5
  assign b_i_k_9_i_j_1 = _T_2599;	// matmul/matmul-hw.mlir:14971:5
  //PROBE: b_i_k_9_i_j_1	// matmul/matmul-hw.mlir:14972:5
  assign c_prev_i_k_9_i_j_1 = C_reg_bank9_p0_rd_data_2427;	// matmul/matmul-hw.mlir:14683:36, :14974:5
  //PROBE: c_prev_i_k_9_i_j_1	// matmul/matmul-hw.mlir:14975:5
  assign tk_i_k_9_i_j_1 = _T_2819;	// matmul/matmul-hw.mlir:14977:5
  //PROBE: tk_i_k_9_i_j_1	// matmul/matmul-hw.mlir:14978:5
  wire [31:0] _T_3027 = mult_inst25_result + C_reg_bank9_p0_rd_data_2427;	// matmul/matmul-hw.mlir:14683:36, :14965:27, :14979:13
  assign c_i_k_9_i_j_1 = _T_3027;	// matmul/matmul-hw.mlir:14981:5
  //PROBE: c_i_k_9_i_j_1	// matmul/matmul-hw.mlir:14982:5
  assign _T_1253 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14983:13
  assign _T_1252 = _T_2863 ? _T_3027 : 32'bx;	// matmul/matmul-hw.mlir:9287:19, :14984:13
  localparam [3:0] _T_3029 = 4'h0;	// matmul/matmul-hw.mlir:14987:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:14988:5
    if (rst)	// matmul/matmul-hw.mlir:14988:5
      i_k_next_3028 <= _T_3029;	// matmul/matmul-hw.mlir:14991:7
    else	// matmul/matmul-hw.mlir:14988:5
      i_k_next_3028 <= i_k_next_3025;	// matmul/matmul-hw.mlir:14956:13, :14989:7
  end // always @(posedge)
  assign _T_1251 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14993:13
  assign _T_1250 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14994:13
  mult mult_inst26 (	// matmul/matmul-hw.mlir:14995:27
    .a      (A_reg_bank26_p0_rd_data),	// matmul/matmul-hw.mlir:12241:32
    .b      (_T_2615),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst26_result)
  );
  assign _T_1249 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :14996:13
  assign a_i_k_10_i_j_1 = A_reg_bank26_p0_rd_data;	// matmul/matmul-hw.mlir:12241:32, :14998:5
  //PROBE: a_i_k_10_i_j_1	// matmul/matmul-hw.mlir:14999:5
  assign b_i_k_10_i_j_1 = _T_2615;	// matmul/matmul-hw.mlir:15001:5
  //PROBE: b_i_k_10_i_j_1	// matmul/matmul-hw.mlir:15002:5
  assign c_prev_i_k_10_i_j_1 = C_reg_bank10_p0_rd_data_2426;	// matmul/matmul-hw.mlir:14684:37, :15004:5
  //PROBE: c_prev_i_k_10_i_j_1	// matmul/matmul-hw.mlir:15005:5
  assign tk_i_k_10_i_j_1 = _T_2830;	// matmul/matmul-hw.mlir:15007:5
  //PROBE: tk_i_k_10_i_j_1	// matmul/matmul-hw.mlir:15008:5
  wire [31:0] _T_3030 = mult_inst26_result + C_reg_bank10_p0_rd_data_2426;	// matmul/matmul-hw.mlir:14684:37, :14995:27, :15009:13
  assign c_i_k_10_i_j_1 = _T_3030;	// matmul/matmul-hw.mlir:15011:5
  //PROBE: c_i_k_10_i_j_1	// matmul/matmul-hw.mlir:15012:5
  assign _T_1248 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15013:13
  assign _T_1247 = _T_2874 ? _T_3030 : 32'bx;	// matmul/matmul-hw.mlir:9282:19, :15014:13
  localparam [3:0] _T_3032 = 4'h0;	// matmul/matmul-hw.mlir:15017:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15018:5
    if (rst)	// matmul/matmul-hw.mlir:15018:5
      i_k_next_3031 <= _T_3032;	// matmul/matmul-hw.mlir:15021:7
    else	// matmul/matmul-hw.mlir:15018:5
      i_k_next_3031 <= i_k_next_3028;	// matmul/matmul-hw.mlir:14986:13, :15019:7
  end // always @(posedge)
  assign _T_1246 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15023:13
  assign _T_1245 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15024:13
  mult mult_inst27 (	// matmul/matmul-hw.mlir:15025:27
    .a      (A_reg_bank27_p0_rd_data),	// matmul/matmul-hw.mlir:12242:32
    .b      (_T_2631),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst27_result)
  );
  assign _T_1244 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15026:13
  assign a_i_k_11_i_j_1 = A_reg_bank27_p0_rd_data;	// matmul/matmul-hw.mlir:12242:32, :15028:5
  //PROBE: a_i_k_11_i_j_1	// matmul/matmul-hw.mlir:15029:5
  assign b_i_k_11_i_j_1 = _T_2631;	// matmul/matmul-hw.mlir:15031:5
  //PROBE: b_i_k_11_i_j_1	// matmul/matmul-hw.mlir:15032:5
  assign c_prev_i_k_11_i_j_1 = C_reg_bank11_p0_rd_data_2425;	// matmul/matmul-hw.mlir:14685:37, :15034:5
  //PROBE: c_prev_i_k_11_i_j_1	// matmul/matmul-hw.mlir:15035:5
  assign tk_i_k_11_i_j_1 = _T_2841;	// matmul/matmul-hw.mlir:15037:5
  //PROBE: tk_i_k_11_i_j_1	// matmul/matmul-hw.mlir:15038:5
  wire [31:0] _T_3033 = mult_inst27_result + C_reg_bank11_p0_rd_data_2425;	// matmul/matmul-hw.mlir:14685:37, :15025:27, :15039:13
  assign c_i_k_11_i_j_1 = _T_3033;	// matmul/matmul-hw.mlir:15041:5
  //PROBE: c_i_k_11_i_j_1	// matmul/matmul-hw.mlir:15042:5
  assign _T_1243 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15043:13
  assign _T_1242 = _T_2885 ? _T_3033 : 32'bx;	// matmul/matmul-hw.mlir:9277:19, :15044:13
  localparam [3:0] _T_3035 = 4'h0;	// matmul/matmul-hw.mlir:15047:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15048:5
    if (rst)	// matmul/matmul-hw.mlir:15048:5
      i_k_next_3034 <= _T_3035;	// matmul/matmul-hw.mlir:15051:7
    else	// matmul/matmul-hw.mlir:15048:5
      i_k_next_3034 <= i_k_next_3031;	// matmul/matmul-hw.mlir:15016:13, :15049:7
  end // always @(posedge)
  assign _T_1241 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15053:13
  assign _T_1240 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15054:13
  mult mult_inst28 (	// matmul/matmul-hw.mlir:15055:27
    .a      (A_reg_bank28_p0_rd_data),	// matmul/matmul-hw.mlir:12243:32
    .b      (_T_2647),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst28_result)
  );
  assign _T_1239 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15056:13
  assign a_i_k_12_i_j_1 = A_reg_bank28_p0_rd_data;	// matmul/matmul-hw.mlir:12243:32, :15058:5
  //PROBE: a_i_k_12_i_j_1	// matmul/matmul-hw.mlir:15059:5
  assign b_i_k_12_i_j_1 = _T_2647;	// matmul/matmul-hw.mlir:15061:5
  //PROBE: b_i_k_12_i_j_1	// matmul/matmul-hw.mlir:15062:5
  assign c_prev_i_k_12_i_j_1 = C_reg_bank12_p0_rd_data_2424;	// matmul/matmul-hw.mlir:14686:37, :15064:5
  //PROBE: c_prev_i_k_12_i_j_1	// matmul/matmul-hw.mlir:15065:5
  assign tk_i_k_12_i_j_1 = _T_2852;	// matmul/matmul-hw.mlir:15067:5
  //PROBE: tk_i_k_12_i_j_1	// matmul/matmul-hw.mlir:15068:5
  wire [31:0] _T_3036 = mult_inst28_result + C_reg_bank12_p0_rd_data_2424;	// matmul/matmul-hw.mlir:14686:37, :15055:27, :15069:13
  assign c_i_k_12_i_j_1 = _T_3036;	// matmul/matmul-hw.mlir:15071:5
  //PROBE: c_i_k_12_i_j_1	// matmul/matmul-hw.mlir:15072:5
  assign _T_1238 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15073:13
  assign _T_1237 = _T_2892 ? _T_3036 : 32'bx;	// matmul/matmul-hw.mlir:9272:19, :15074:13
  localparam [3:0] _T_3038 = 4'h0;	// matmul/matmul-hw.mlir:15077:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15078:5
    if (rst)	// matmul/matmul-hw.mlir:15078:5
      i_k_next_3037 <= _T_3038;	// matmul/matmul-hw.mlir:15081:7
    else	// matmul/matmul-hw.mlir:15078:5
      i_k_next_3037 <= i_k_next_3034;	// matmul/matmul-hw.mlir:15046:13, :15079:7
  end // always @(posedge)
  assign _T_1236 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15083:13
  assign _T_1235 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15084:13
  mult mult_inst29 (	// matmul/matmul-hw.mlir:15085:27
    .a      (A_reg_bank29_p0_rd_data),	// matmul/matmul-hw.mlir:12244:32
    .b      (_T_2663),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst29_result)
  );
  assign _T_1234 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15086:13
  assign a_i_k_13_i_j_1 = A_reg_bank29_p0_rd_data;	// matmul/matmul-hw.mlir:12244:32, :15088:5
  //PROBE: a_i_k_13_i_j_1	// matmul/matmul-hw.mlir:15089:5
  assign b_i_k_13_i_j_1 = _T_2663;	// matmul/matmul-hw.mlir:15091:5
  //PROBE: b_i_k_13_i_j_1	// matmul/matmul-hw.mlir:15092:5
  assign c_prev_i_k_13_i_j_1 = C_reg_bank13_p0_rd_data_2423;	// matmul/matmul-hw.mlir:14687:37, :15094:5
  //PROBE: c_prev_i_k_13_i_j_1	// matmul/matmul-hw.mlir:15095:5
  assign tk_i_k_13_i_j_1 = _T_2863;	// matmul/matmul-hw.mlir:15097:5
  //PROBE: tk_i_k_13_i_j_1	// matmul/matmul-hw.mlir:15098:5
  wire [31:0] _T_3039 = mult_inst29_result + C_reg_bank13_p0_rd_data_2423;	// matmul/matmul-hw.mlir:14687:37, :15085:27, :15099:13
  assign c_i_k_13_i_j_1 = _T_3039;	// matmul/matmul-hw.mlir:15101:5
  //PROBE: c_i_k_13_i_j_1	// matmul/matmul-hw.mlir:15102:5
  assign _T_1233 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15103:13
  assign _T_1232 = _T_2897 ? _T_3039 : 32'bx;	// matmul/matmul-hw.mlir:9267:19, :15104:13
  localparam [3:0] _T_3041 = 4'h0;	// matmul/matmul-hw.mlir:15107:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15108:5
    if (rst)	// matmul/matmul-hw.mlir:15108:5
      i_k_next_3040 <= _T_3041;	// matmul/matmul-hw.mlir:15111:7
    else	// matmul/matmul-hw.mlir:15108:5
      i_k_next_3040 <= i_k_next_3037;	// matmul/matmul-hw.mlir:15076:13, :15109:7
  end // always @(posedge)
  assign _T_1231 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15113:13
  assign _T_1230 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15114:13
  mult mult_inst30 (	// matmul/matmul-hw.mlir:15115:27
    .a      (A_reg_bank30_p0_rd_data),	// matmul/matmul-hw.mlir:12245:32
    .b      (_T_2679),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst30_result)
  );
  assign _T_1229 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15116:13
  assign a_i_k_14_i_j_1 = A_reg_bank30_p0_rd_data;	// matmul/matmul-hw.mlir:12245:32, :15118:5
  //PROBE: a_i_k_14_i_j_1	// matmul/matmul-hw.mlir:15119:5
  assign b_i_k_14_i_j_1 = _T_2679;	// matmul/matmul-hw.mlir:15121:5
  //PROBE: b_i_k_14_i_j_1	// matmul/matmul-hw.mlir:15122:5
  assign c_prev_i_k_14_i_j_1 = C_reg_bank14_p0_rd_data_2422;	// matmul/matmul-hw.mlir:14688:37, :15124:5
  //PROBE: c_prev_i_k_14_i_j_1	// matmul/matmul-hw.mlir:15125:5
  assign tk_i_k_14_i_j_1 = _T_2874;	// matmul/matmul-hw.mlir:15127:5
  //PROBE: tk_i_k_14_i_j_1	// matmul/matmul-hw.mlir:15128:5
  wire [31:0] _T_3042 = mult_inst30_result + C_reg_bank14_p0_rd_data_2422;	// matmul/matmul-hw.mlir:14688:37, :15115:27, :15129:13
  assign c_i_k_14_i_j_1 = _T_3042;	// matmul/matmul-hw.mlir:15131:5
  //PROBE: c_i_k_14_i_j_1	// matmul/matmul-hw.mlir:15132:5
  assign _T_1228 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15133:13
  assign _T_1227 = _T_2902 ? _T_3042 : 32'bx;	// matmul/matmul-hw.mlir:9262:19, :15134:13
  localparam [3:0] _T_3044 = 4'h0;	// matmul/matmul-hw.mlir:15137:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15138:5
    if (rst)	// matmul/matmul-hw.mlir:15138:5
      i_k_next_3043 <= _T_3044;	// matmul/matmul-hw.mlir:15141:7
    else	// matmul/matmul-hw.mlir:15138:5
      i_k_next_3043 <= i_k_next_3040;	// matmul/matmul-hw.mlir:15106:13, :15139:7
  end // always @(posedge)
  assign _T_1226 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15143:13
  assign _T_1225 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15144:13
  mult mult_inst31 (	// matmul/matmul-hw.mlir:15145:27
    .a      (A_reg_bank31_p0_rd_data),	// matmul/matmul-hw.mlir:12246:32
    .b      (_T_2695),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst31_result)
  );
  assign _T_1224 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15146:13
  assign a_i_k_15_i_j_1 = A_reg_bank31_p0_rd_data;	// matmul/matmul-hw.mlir:12246:32, :15148:5
  //PROBE: a_i_k_15_i_j_1	// matmul/matmul-hw.mlir:15149:5
  assign b_i_k_15_i_j_1 = _T_2695;	// matmul/matmul-hw.mlir:15151:5
  //PROBE: b_i_k_15_i_j_1	// matmul/matmul-hw.mlir:15152:5
  assign c_prev_i_k_15_i_j_1 = C_reg_bank15_p0_rd_data_2421;	// matmul/matmul-hw.mlir:14689:37, :15154:5
  //PROBE: c_prev_i_k_15_i_j_1	// matmul/matmul-hw.mlir:15155:5
  assign tk_i_k_15_i_j_1 = _T_2885;	// matmul/matmul-hw.mlir:15157:5
  //PROBE: tk_i_k_15_i_j_1	// matmul/matmul-hw.mlir:15158:5
  wire [31:0] _T_3045 = mult_inst31_result + C_reg_bank15_p0_rd_data_2421;	// matmul/matmul-hw.mlir:14689:37, :15145:27, :15159:13
  assign c_i_k_15_i_j_1 = _T_3045;	// matmul/matmul-hw.mlir:15161:5
  //PROBE: c_i_k_15_i_j_1	// matmul/matmul-hw.mlir:15162:5
  assign _T_1223 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15163:13
  assign _T_1222 = _T_2907 ? _T_3045 : 32'bx;	// matmul/matmul-hw.mlir:9257:19, :15164:13
  localparam [3:0] _T_3047 = 4'h0;	// matmul/matmul-hw.mlir:15167:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15168:5
    if (rst)	// matmul/matmul-hw.mlir:15168:5
      i_k_next_3046 <= _T_3047;	// matmul/matmul-hw.mlir:15171:7
    else	// matmul/matmul-hw.mlir:15168:5
      i_k_next_3046 <= i_k_next_3043;	// matmul/matmul-hw.mlir:15136:13, :15169:7
  end // always @(posedge)
  assign _T_1221 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15173:13
  wire [3:0][3:0] _T_3049 = i_delayed_3048;	// matmul/matmul-hw.mlir:15175:13
  wire [3:0][3:0] _T_3050 = {_T_3049[2'h0+:3], {{i_k_next_3046}}};	// matmul/matmul-hw.mlir:15166:13, :15176:19, :15177:13, :15178:13, :15179:13
  wire [3:0][3:0] _T_3051 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:15180:19, :15181:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15182:5
    if (rst)	// matmul/matmul-hw.mlir:15182:5
      i_delayed_3048 <= _T_3051;	// matmul/matmul-hw.mlir:15185:7
    else	// matmul/matmul-hw.mlir:15182:5
      i_delayed_3048 <= _T_3050;	// matmul/matmul-hw.mlir:15183:7
  end // always @(posedge)
  assign _T_1220 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15189:13
  assign _T_1219 = _T_2912 ? i_delayed_3048[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:9254:18, :15175:13, :15187:20, :15188:13, :15190:13
  assign _T_1218 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15191:13
  assign _T_1217 = _T_2912 ? C_reg_bank16_p0_rd_data_2420 : 32'bx;	// matmul/matmul-hw.mlir:9252:19, :14690:37, :15192:13
  localparam [3:0] _T_3053 = 4'h0;	// matmul/matmul-hw.mlir:15195:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15196:5
    if (rst)	// matmul/matmul-hw.mlir:15196:5
      i_j_next_3052 <= _T_3053;	// matmul/matmul-hw.mlir:15199:7
    else	// matmul/matmul-hw.mlir:15196:5
      i_j_next_3052 <= i_j_next;	// matmul/matmul-hw.mlir:14599:13, :15197:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3054 (	// matmul/matmul-hw.mlir:15269:36
    .p0_rd_en   (_T_1212),	// matmul/matmul-hw.mlir:15291:13
    .p1_wr_en   (_T_1216),	// matmul/matmul-hw.mlir:15286:13
    .p1_wr_data (_T_1215),	// matmul/matmul-hw.mlir:15287:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2419)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3055 (	// matmul/matmul-hw.mlir:15270:36
    .p0_rd_en   (_T_1207),	// matmul/matmul-hw.mlir:15321:13
    .p1_wr_en   (_T_1211),	// matmul/matmul-hw.mlir:15308:13
    .p1_wr_data (_T_1210),	// matmul/matmul-hw.mlir:15309:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2418)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3056 (	// matmul/matmul-hw.mlir:15271:36
    .p0_rd_en   (_T_1202),	// matmul/matmul-hw.mlir:15351:13
    .p1_wr_en   (_T_1206),	// matmul/matmul-hw.mlir:15338:13
    .p1_wr_data (_T_1205),	// matmul/matmul-hw.mlir:15339:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2417)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3057 (	// matmul/matmul-hw.mlir:15272:36
    .p0_rd_en   (_T_1197),	// matmul/matmul-hw.mlir:15381:13
    .p1_wr_en   (_T_1201),	// matmul/matmul-hw.mlir:15368:13
    .p1_wr_data (_T_1200),	// matmul/matmul-hw.mlir:15369:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2416)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3058 (	// matmul/matmul-hw.mlir:15273:36
    .p0_rd_en   (_T_1192),	// matmul/matmul-hw.mlir:15411:13
    .p1_wr_en   (_T_1196),	// matmul/matmul-hw.mlir:15398:13
    .p1_wr_data (_T_1195),	// matmul/matmul-hw.mlir:15399:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2415)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3059 (	// matmul/matmul-hw.mlir:15274:36
    .p0_rd_en   (_T_1187),	// matmul/matmul-hw.mlir:15441:13
    .p1_wr_en   (_T_1191),	// matmul/matmul-hw.mlir:15428:13
    .p1_wr_data (_T_1190),	// matmul/matmul-hw.mlir:15429:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2414)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3060 (	// matmul/matmul-hw.mlir:15275:36
    .p0_rd_en   (_T_1182),	// matmul/matmul-hw.mlir:15471:13
    .p1_wr_en   (_T_1186),	// matmul/matmul-hw.mlir:15458:13
    .p1_wr_data (_T_1185),	// matmul/matmul-hw.mlir:15459:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2413)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3061 (	// matmul/matmul-hw.mlir:15276:36
    .p0_rd_en   (_T_1177),	// matmul/matmul-hw.mlir:15501:13
    .p1_wr_en   (_T_1181),	// matmul/matmul-hw.mlir:15488:13
    .p1_wr_data (_T_1180),	// matmul/matmul-hw.mlir:15489:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2412)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3062 (	// matmul/matmul-hw.mlir:15277:36
    .p0_rd_en   (_T_1172),	// matmul/matmul-hw.mlir:15531:13
    .p1_wr_en   (_T_1176),	// matmul/matmul-hw.mlir:15518:13
    .p1_wr_data (_T_1175),	// matmul/matmul-hw.mlir:15519:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2411)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3063 (	// matmul/matmul-hw.mlir:15278:36
    .p0_rd_en   (_T_1167),	// matmul/matmul-hw.mlir:15561:13
    .p1_wr_en   (_T_1171),	// matmul/matmul-hw.mlir:15548:13
    .p1_wr_data (_T_1170),	// matmul/matmul-hw.mlir:15549:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2410)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3064 (	// matmul/matmul-hw.mlir:15279:37
    .p0_rd_en   (_T_1162),	// matmul/matmul-hw.mlir:15591:13
    .p1_wr_en   (_T_1166),	// matmul/matmul-hw.mlir:15578:13
    .p1_wr_data (_T_1165),	// matmul/matmul-hw.mlir:15579:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2409)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3065 (	// matmul/matmul-hw.mlir:15280:37
    .p0_rd_en   (_T_1157),	// matmul/matmul-hw.mlir:15621:13
    .p1_wr_en   (_T_1161),	// matmul/matmul-hw.mlir:15608:13
    .p1_wr_data (_T_1160),	// matmul/matmul-hw.mlir:15609:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2408)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3066 (	// matmul/matmul-hw.mlir:15281:37
    .p0_rd_en   (_T_1152),	// matmul/matmul-hw.mlir:15651:13
    .p1_wr_en   (_T_1156),	// matmul/matmul-hw.mlir:15638:13
    .p1_wr_data (_T_1155),	// matmul/matmul-hw.mlir:15639:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2407)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3067 (	// matmul/matmul-hw.mlir:15282:37
    .p0_rd_en   (_T_1147),	// matmul/matmul-hw.mlir:15681:13
    .p1_wr_en   (_T_1151),	// matmul/matmul-hw.mlir:15668:13
    .p1_wr_data (_T_1150),	// matmul/matmul-hw.mlir:15669:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2406)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3068 (	// matmul/matmul-hw.mlir:15283:37
    .p0_rd_en   (_T_1142),	// matmul/matmul-hw.mlir:15711:13
    .p1_wr_en   (_T_1146),	// matmul/matmul-hw.mlir:15698:13
    .p1_wr_data (_T_1145),	// matmul/matmul-hw.mlir:15699:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2405)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3069 (	// matmul/matmul-hw.mlir:15284:37
    .p0_rd_en   (_T_1137),	// matmul/matmul-hw.mlir:15741:13
    .p1_wr_en   (_T_1141),	// matmul/matmul-hw.mlir:15728:13
    .p1_wr_data (_T_1140),	// matmul/matmul-hw.mlir:15729:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2404)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3070 (	// matmul/matmul-hw.mlir:15285:37
    .p0_rd_en   (_T_1134),	// matmul/matmul-hw.mlir:15768:13
    .p1_wr_en   (_T_1136),	// matmul/matmul-hw.mlir:15758:13
    .p1_wr_data (_T_1135),	// matmul/matmul-hw.mlir:15759:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2403)
  );
  assign _T_1216 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15286:13
  assign _T_1215 = _T_2764 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :9250:19, :15287:13
  assign _T_1214 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15288:13
  assign _T_1213 = _T_2753 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15289:13
  mult mult_inst32 (	// matmul/matmul-hw.mlir:15290:27
    .a      (A_reg_bank32_p0_rd_data),	// matmul/matmul-hw.mlir:12247:32
    .b      (_T_2456),
    .t      (_T_2753),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst32_result)
  );
  assign _T_1212 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15291:13
  assign a_i_k_0_i_j_2 = A_reg_bank32_p0_rd_data;	// matmul/matmul-hw.mlir:12247:32, :15293:5
  //PROBE: a_i_k_0_i_j_2	// matmul/matmul-hw.mlir:15294:5
  assign b_i_k_0_i_j_2 = _T_2456;	// matmul/matmul-hw.mlir:15296:5
  //PROBE: b_i_k_0_i_j_2	// matmul/matmul-hw.mlir:15297:5
  assign c_prev_i_k_0_i_j_2 = C_reg_bank0_p0_rd_data_2419;	// matmul/matmul-hw.mlir:15269:36, :15299:5
  //PROBE: c_prev_i_k_0_i_j_2	// matmul/matmul-hw.mlir:15300:5
  assign tk_i_k_0_i_j_2 = _T_2731;	// matmul/matmul-hw.mlir:15302:5
  //PROBE: tk_i_k_0_i_j_2	// matmul/matmul-hw.mlir:15303:5
  wire [31:0] _T_3071 = mult_inst32_result + C_reg_bank0_p0_rd_data_2419;	// matmul/matmul-hw.mlir:15269:36, :15290:27, :15304:13
  assign c_i_k_0_i_j_2 = _T_3071;	// matmul/matmul-hw.mlir:15306:5
  //PROBE: c_i_k_0_i_j_2	// matmul/matmul-hw.mlir:15307:5
  assign _T_1211 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15308:13
  assign _T_1210 = _T_2775 ? _T_3071 : 32'bx;	// matmul/matmul-hw.mlir:9245:19, :15309:13
  localparam [3:0] _T_3073 = 4'h0;	// matmul/matmul-hw.mlir:15312:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15313:5
    if (rst)	// matmul/matmul-hw.mlir:15313:5
      i_k_next_3072 <= _T_3073;	// matmul/matmul-hw.mlir:15316:7
    else	// matmul/matmul-hw.mlir:15313:5
      i_k_next_3072 <= i_j_next_3052;	// matmul/matmul-hw.mlir:15194:13, :15314:7
  end // always @(posedge)
  assign _T_1209 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15318:13
  assign _T_1208 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15319:13
  mult mult_inst33 (	// matmul/matmul-hw.mlir:15320:27
    .a      (A_reg_bank33_p0_rd_data),	// matmul/matmul-hw.mlir:12248:32
    .b      (_T_2472),
    .t      (_T_2764),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst33_result)
  );
  assign _T_1207 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15321:13
  assign a_i_k_1_i_j_2 = A_reg_bank33_p0_rd_data;	// matmul/matmul-hw.mlir:12248:32, :15323:5
  //PROBE: a_i_k_1_i_j_2	// matmul/matmul-hw.mlir:15324:5
  assign b_i_k_1_i_j_2 = _T_2472;	// matmul/matmul-hw.mlir:15326:5
  //PROBE: b_i_k_1_i_j_2	// matmul/matmul-hw.mlir:15327:5
  assign c_prev_i_k_1_i_j_2 = C_reg_bank1_p0_rd_data_2418;	// matmul/matmul-hw.mlir:15270:36, :15329:5
  //PROBE: c_prev_i_k_1_i_j_2	// matmul/matmul-hw.mlir:15330:5
  assign tk_i_k_1_i_j_2 = _T_2742;	// matmul/matmul-hw.mlir:15332:5
  //PROBE: tk_i_k_1_i_j_2	// matmul/matmul-hw.mlir:15333:5
  wire [31:0] _T_3074 = mult_inst33_result + C_reg_bank1_p0_rd_data_2418;	// matmul/matmul-hw.mlir:15270:36, :15320:27, :15334:13
  assign c_i_k_1_i_j_2 = _T_3074;	// matmul/matmul-hw.mlir:15336:5
  //PROBE: c_i_k_1_i_j_2	// matmul/matmul-hw.mlir:15337:5
  assign _T_1206 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15338:13
  assign _T_1205 = _T_2786 ? _T_3074 : 32'bx;	// matmul/matmul-hw.mlir:9240:19, :15339:13
  localparam [3:0] _T_3076 = 4'h0;	// matmul/matmul-hw.mlir:15342:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15343:5
    if (rst)	// matmul/matmul-hw.mlir:15343:5
      i_k_next_3075 <= _T_3076;	// matmul/matmul-hw.mlir:15346:7
    else	// matmul/matmul-hw.mlir:15343:5
      i_k_next_3075 <= i_k_next_3072;	// matmul/matmul-hw.mlir:15311:13, :15344:7
  end // always @(posedge)
  assign _T_1204 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15348:13
  assign _T_1203 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15349:13
  mult mult_inst34 (	// matmul/matmul-hw.mlir:15350:27
    .a      (A_reg_bank34_p0_rd_data),	// matmul/matmul-hw.mlir:12249:32
    .b      (_T_2488),
    .t      (_T_2775),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst34_result)
  );
  assign _T_1202 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15351:13
  assign a_i_k_2_i_j_2 = A_reg_bank34_p0_rd_data;	// matmul/matmul-hw.mlir:12249:32, :15353:5
  //PROBE: a_i_k_2_i_j_2	// matmul/matmul-hw.mlir:15354:5
  assign b_i_k_2_i_j_2 = _T_2488;	// matmul/matmul-hw.mlir:15356:5
  //PROBE: b_i_k_2_i_j_2	// matmul/matmul-hw.mlir:15357:5
  assign c_prev_i_k_2_i_j_2 = C_reg_bank2_p0_rd_data_2417;	// matmul/matmul-hw.mlir:15271:36, :15359:5
  //PROBE: c_prev_i_k_2_i_j_2	// matmul/matmul-hw.mlir:15360:5
  assign tk_i_k_2_i_j_2 = _T_2753;	// matmul/matmul-hw.mlir:15362:5
  //PROBE: tk_i_k_2_i_j_2	// matmul/matmul-hw.mlir:15363:5
  wire [31:0] _T_3077 = mult_inst34_result + C_reg_bank2_p0_rd_data_2417;	// matmul/matmul-hw.mlir:15271:36, :15350:27, :15364:13
  assign c_i_k_2_i_j_2 = _T_3077;	// matmul/matmul-hw.mlir:15366:5
  //PROBE: c_i_k_2_i_j_2	// matmul/matmul-hw.mlir:15367:5
  assign _T_1201 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15368:13
  assign _T_1200 = _T_2797 ? _T_3077 : 32'bx;	// matmul/matmul-hw.mlir:9235:19, :15369:13
  localparam [3:0] _T_3079 = 4'h0;	// matmul/matmul-hw.mlir:15372:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15373:5
    if (rst)	// matmul/matmul-hw.mlir:15373:5
      i_k_next_3078 <= _T_3079;	// matmul/matmul-hw.mlir:15376:7
    else	// matmul/matmul-hw.mlir:15373:5
      i_k_next_3078 <= i_k_next_3075;	// matmul/matmul-hw.mlir:15341:13, :15374:7
  end // always @(posedge)
  assign _T_1199 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15378:13
  assign _T_1198 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15379:13
  mult mult_inst35 (	// matmul/matmul-hw.mlir:15380:27
    .a      (A_reg_bank35_p0_rd_data),	// matmul/matmul-hw.mlir:12250:32
    .b      (_T_2504),
    .t      (_T_2786),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst35_result)
  );
  assign _T_1197 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15381:13
  assign a_i_k_3_i_j_2 = A_reg_bank35_p0_rd_data;	// matmul/matmul-hw.mlir:12250:32, :15383:5
  //PROBE: a_i_k_3_i_j_2	// matmul/matmul-hw.mlir:15384:5
  assign b_i_k_3_i_j_2 = _T_2504;	// matmul/matmul-hw.mlir:15386:5
  //PROBE: b_i_k_3_i_j_2	// matmul/matmul-hw.mlir:15387:5
  assign c_prev_i_k_3_i_j_2 = C_reg_bank3_p0_rd_data_2416;	// matmul/matmul-hw.mlir:15272:36, :15389:5
  //PROBE: c_prev_i_k_3_i_j_2	// matmul/matmul-hw.mlir:15390:5
  assign tk_i_k_3_i_j_2 = _T_2764;	// matmul/matmul-hw.mlir:15392:5
  //PROBE: tk_i_k_3_i_j_2	// matmul/matmul-hw.mlir:15393:5
  wire [31:0] _T_3080 = mult_inst35_result + C_reg_bank3_p0_rd_data_2416;	// matmul/matmul-hw.mlir:15272:36, :15380:27, :15394:13
  assign c_i_k_3_i_j_2 = _T_3080;	// matmul/matmul-hw.mlir:15396:5
  //PROBE: c_i_k_3_i_j_2	// matmul/matmul-hw.mlir:15397:5
  assign _T_1196 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15398:13
  assign _T_1195 = _T_2808 ? _T_3080 : 32'bx;	// matmul/matmul-hw.mlir:9230:19, :15399:13
  localparam [3:0] _T_3082 = 4'h0;	// matmul/matmul-hw.mlir:15402:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15403:5
    if (rst)	// matmul/matmul-hw.mlir:15403:5
      i_k_next_3081 <= _T_3082;	// matmul/matmul-hw.mlir:15406:7
    else	// matmul/matmul-hw.mlir:15403:5
      i_k_next_3081 <= i_k_next_3078;	// matmul/matmul-hw.mlir:15371:13, :15404:7
  end // always @(posedge)
  assign _T_1194 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15408:13
  assign _T_1193 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15409:13
  mult mult_inst36 (	// matmul/matmul-hw.mlir:15410:27
    .a      (A_reg_bank36_p0_rd_data),	// matmul/matmul-hw.mlir:12251:32
    .b      (_T_2520),
    .t      (_T_2797),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst36_result)
  );
  assign _T_1192 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15411:13
  assign a_i_k_4_i_j_2 = A_reg_bank36_p0_rd_data;	// matmul/matmul-hw.mlir:12251:32, :15413:5
  //PROBE: a_i_k_4_i_j_2	// matmul/matmul-hw.mlir:15414:5
  assign b_i_k_4_i_j_2 = _T_2520;	// matmul/matmul-hw.mlir:15416:5
  //PROBE: b_i_k_4_i_j_2	// matmul/matmul-hw.mlir:15417:5
  assign c_prev_i_k_4_i_j_2 = C_reg_bank4_p0_rd_data_2415;	// matmul/matmul-hw.mlir:15273:36, :15419:5
  //PROBE: c_prev_i_k_4_i_j_2	// matmul/matmul-hw.mlir:15420:5
  assign tk_i_k_4_i_j_2 = _T_2775;	// matmul/matmul-hw.mlir:15422:5
  //PROBE: tk_i_k_4_i_j_2	// matmul/matmul-hw.mlir:15423:5
  wire [31:0] _T_3083 = mult_inst36_result + C_reg_bank4_p0_rd_data_2415;	// matmul/matmul-hw.mlir:15273:36, :15410:27, :15424:13
  assign c_i_k_4_i_j_2 = _T_3083;	// matmul/matmul-hw.mlir:15426:5
  //PROBE: c_i_k_4_i_j_2	// matmul/matmul-hw.mlir:15427:5
  assign _T_1191 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15428:13
  assign _T_1190 = _T_2819 ? _T_3083 : 32'bx;	// matmul/matmul-hw.mlir:9225:19, :15429:13
  localparam [3:0] _T_3085 = 4'h0;	// matmul/matmul-hw.mlir:15432:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15433:5
    if (rst)	// matmul/matmul-hw.mlir:15433:5
      i_k_next_3084 <= _T_3085;	// matmul/matmul-hw.mlir:15436:7
    else	// matmul/matmul-hw.mlir:15433:5
      i_k_next_3084 <= i_k_next_3081;	// matmul/matmul-hw.mlir:15401:13, :15434:7
  end // always @(posedge)
  assign _T_1189 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15438:13
  assign _T_1188 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15439:13
  mult mult_inst37 (	// matmul/matmul-hw.mlir:15440:27
    .a      (A_reg_bank37_p0_rd_data),	// matmul/matmul-hw.mlir:12252:32
    .b      (_T_2536),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst37_result)
  );
  assign _T_1187 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15441:13
  assign a_i_k_5_i_j_2 = A_reg_bank37_p0_rd_data;	// matmul/matmul-hw.mlir:12252:32, :15443:5
  //PROBE: a_i_k_5_i_j_2	// matmul/matmul-hw.mlir:15444:5
  assign b_i_k_5_i_j_2 = _T_2536;	// matmul/matmul-hw.mlir:15446:5
  //PROBE: b_i_k_5_i_j_2	// matmul/matmul-hw.mlir:15447:5
  assign c_prev_i_k_5_i_j_2 = C_reg_bank5_p0_rd_data_2414;	// matmul/matmul-hw.mlir:15274:36, :15449:5
  //PROBE: c_prev_i_k_5_i_j_2	// matmul/matmul-hw.mlir:15450:5
  assign tk_i_k_5_i_j_2 = _T_2786;	// matmul/matmul-hw.mlir:15452:5
  //PROBE: tk_i_k_5_i_j_2	// matmul/matmul-hw.mlir:15453:5
  wire [31:0] _T_3086 = mult_inst37_result + C_reg_bank5_p0_rd_data_2414;	// matmul/matmul-hw.mlir:15274:36, :15440:27, :15454:13
  assign c_i_k_5_i_j_2 = _T_3086;	// matmul/matmul-hw.mlir:15456:5
  //PROBE: c_i_k_5_i_j_2	// matmul/matmul-hw.mlir:15457:5
  assign _T_1186 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15458:13
  assign _T_1185 = _T_2830 ? _T_3086 : 32'bx;	// matmul/matmul-hw.mlir:9220:19, :15459:13
  localparam [3:0] _T_3088 = 4'h0;	// matmul/matmul-hw.mlir:15462:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15463:5
    if (rst)	// matmul/matmul-hw.mlir:15463:5
      i_k_next_3087 <= _T_3088;	// matmul/matmul-hw.mlir:15466:7
    else	// matmul/matmul-hw.mlir:15463:5
      i_k_next_3087 <= i_k_next_3084;	// matmul/matmul-hw.mlir:15431:13, :15464:7
  end // always @(posedge)
  assign _T_1184 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15468:13
  assign _T_1183 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15469:13
  mult mult_inst38 (	// matmul/matmul-hw.mlir:15470:27
    .a      (A_reg_bank38_p0_rd_data),	// matmul/matmul-hw.mlir:12253:32
    .b      (_T_2552),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst38_result)
  );
  assign _T_1182 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15471:13
  assign a_i_k_6_i_j_2 = A_reg_bank38_p0_rd_data;	// matmul/matmul-hw.mlir:12253:32, :15473:5
  //PROBE: a_i_k_6_i_j_2	// matmul/matmul-hw.mlir:15474:5
  assign b_i_k_6_i_j_2 = _T_2552;	// matmul/matmul-hw.mlir:15476:5
  //PROBE: b_i_k_6_i_j_2	// matmul/matmul-hw.mlir:15477:5
  assign c_prev_i_k_6_i_j_2 = C_reg_bank6_p0_rd_data_2413;	// matmul/matmul-hw.mlir:15275:36, :15479:5
  //PROBE: c_prev_i_k_6_i_j_2	// matmul/matmul-hw.mlir:15480:5
  assign tk_i_k_6_i_j_2 = _T_2797;	// matmul/matmul-hw.mlir:15482:5
  //PROBE: tk_i_k_6_i_j_2	// matmul/matmul-hw.mlir:15483:5
  wire [31:0] _T_3089 = mult_inst38_result + C_reg_bank6_p0_rd_data_2413;	// matmul/matmul-hw.mlir:15275:36, :15470:27, :15484:13
  assign c_i_k_6_i_j_2 = _T_3089;	// matmul/matmul-hw.mlir:15486:5
  //PROBE: c_i_k_6_i_j_2	// matmul/matmul-hw.mlir:15487:5
  assign _T_1181 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15488:13
  assign _T_1180 = _T_2841 ? _T_3089 : 32'bx;	// matmul/matmul-hw.mlir:9215:19, :15489:13
  localparam [3:0] _T_3091 = 4'h0;	// matmul/matmul-hw.mlir:15492:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15493:5
    if (rst)	// matmul/matmul-hw.mlir:15493:5
      i_k_next_3090 <= _T_3091;	// matmul/matmul-hw.mlir:15496:7
    else	// matmul/matmul-hw.mlir:15493:5
      i_k_next_3090 <= i_k_next_3087;	// matmul/matmul-hw.mlir:15461:13, :15494:7
  end // always @(posedge)
  assign _T_1179 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15498:13
  assign _T_1178 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15499:13
  mult mult_inst39 (	// matmul/matmul-hw.mlir:15500:27
    .a      (A_reg_bank39_p0_rd_data),	// matmul/matmul-hw.mlir:12254:32
    .b      (_T_2568),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst39_result)
  );
  assign _T_1177 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15501:13
  assign a_i_k_7_i_j_2 = A_reg_bank39_p0_rd_data;	// matmul/matmul-hw.mlir:12254:32, :15503:5
  //PROBE: a_i_k_7_i_j_2	// matmul/matmul-hw.mlir:15504:5
  assign b_i_k_7_i_j_2 = _T_2568;	// matmul/matmul-hw.mlir:15506:5
  //PROBE: b_i_k_7_i_j_2	// matmul/matmul-hw.mlir:15507:5
  assign c_prev_i_k_7_i_j_2 = C_reg_bank7_p0_rd_data_2412;	// matmul/matmul-hw.mlir:15276:36, :15509:5
  //PROBE: c_prev_i_k_7_i_j_2	// matmul/matmul-hw.mlir:15510:5
  assign tk_i_k_7_i_j_2 = _T_2808;	// matmul/matmul-hw.mlir:15512:5
  //PROBE: tk_i_k_7_i_j_2	// matmul/matmul-hw.mlir:15513:5
  wire [31:0] _T_3092 = mult_inst39_result + C_reg_bank7_p0_rd_data_2412;	// matmul/matmul-hw.mlir:15276:36, :15500:27, :15514:13
  assign c_i_k_7_i_j_2 = _T_3092;	// matmul/matmul-hw.mlir:15516:5
  //PROBE: c_i_k_7_i_j_2	// matmul/matmul-hw.mlir:15517:5
  assign _T_1176 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15518:13
  assign _T_1175 = _T_2852 ? _T_3092 : 32'bx;	// matmul/matmul-hw.mlir:9210:19, :15519:13
  localparam [3:0] _T_3094 = 4'h0;	// matmul/matmul-hw.mlir:15522:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15523:5
    if (rst)	// matmul/matmul-hw.mlir:15523:5
      i_k_next_3093 <= _T_3094;	// matmul/matmul-hw.mlir:15526:7
    else	// matmul/matmul-hw.mlir:15523:5
      i_k_next_3093 <= i_k_next_3090;	// matmul/matmul-hw.mlir:15491:13, :15524:7
  end // always @(posedge)
  assign _T_1174 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15528:13
  assign _T_1173 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15529:13
  mult mult_inst40 (	// matmul/matmul-hw.mlir:15530:27
    .a      (A_reg_bank40_p0_rd_data),	// matmul/matmul-hw.mlir:12255:32
    .b      (_T_2584),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst40_result)
  );
  assign _T_1172 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15531:13
  assign a_i_k_8_i_j_2 = A_reg_bank40_p0_rd_data;	// matmul/matmul-hw.mlir:12255:32, :15533:5
  //PROBE: a_i_k_8_i_j_2	// matmul/matmul-hw.mlir:15534:5
  assign b_i_k_8_i_j_2 = _T_2584;	// matmul/matmul-hw.mlir:15536:5
  //PROBE: b_i_k_8_i_j_2	// matmul/matmul-hw.mlir:15537:5
  assign c_prev_i_k_8_i_j_2 = C_reg_bank8_p0_rd_data_2411;	// matmul/matmul-hw.mlir:15277:36, :15539:5
  //PROBE: c_prev_i_k_8_i_j_2	// matmul/matmul-hw.mlir:15540:5
  assign tk_i_k_8_i_j_2 = _T_2819;	// matmul/matmul-hw.mlir:15542:5
  //PROBE: tk_i_k_8_i_j_2	// matmul/matmul-hw.mlir:15543:5
  wire [31:0] _T_3095 = mult_inst40_result + C_reg_bank8_p0_rd_data_2411;	// matmul/matmul-hw.mlir:15277:36, :15530:27, :15544:13
  assign c_i_k_8_i_j_2 = _T_3095;	// matmul/matmul-hw.mlir:15546:5
  //PROBE: c_i_k_8_i_j_2	// matmul/matmul-hw.mlir:15547:5
  assign _T_1171 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15548:13
  assign _T_1170 = _T_2863 ? _T_3095 : 32'bx;	// matmul/matmul-hw.mlir:9205:19, :15549:13
  localparam [3:0] _T_3097 = 4'h0;	// matmul/matmul-hw.mlir:15552:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15553:5
    if (rst)	// matmul/matmul-hw.mlir:15553:5
      i_k_next_3096 <= _T_3097;	// matmul/matmul-hw.mlir:15556:7
    else	// matmul/matmul-hw.mlir:15553:5
      i_k_next_3096 <= i_k_next_3093;	// matmul/matmul-hw.mlir:15521:13, :15554:7
  end // always @(posedge)
  assign _T_1169 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15558:13
  assign _T_1168 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15559:13
  mult mult_inst41 (	// matmul/matmul-hw.mlir:15560:27
    .a      (A_reg_bank41_p0_rd_data),	// matmul/matmul-hw.mlir:12256:32
    .b      (_T_2600),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst41_result)
  );
  assign _T_1167 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15561:13
  assign a_i_k_9_i_j_2 = A_reg_bank41_p0_rd_data;	// matmul/matmul-hw.mlir:12256:32, :15563:5
  //PROBE: a_i_k_9_i_j_2	// matmul/matmul-hw.mlir:15564:5
  assign b_i_k_9_i_j_2 = _T_2600;	// matmul/matmul-hw.mlir:15566:5
  //PROBE: b_i_k_9_i_j_2	// matmul/matmul-hw.mlir:15567:5
  assign c_prev_i_k_9_i_j_2 = C_reg_bank9_p0_rd_data_2410;	// matmul/matmul-hw.mlir:15278:36, :15569:5
  //PROBE: c_prev_i_k_9_i_j_2	// matmul/matmul-hw.mlir:15570:5
  assign tk_i_k_9_i_j_2 = _T_2830;	// matmul/matmul-hw.mlir:15572:5
  //PROBE: tk_i_k_9_i_j_2	// matmul/matmul-hw.mlir:15573:5
  wire [31:0] _T_3098 = mult_inst41_result + C_reg_bank9_p0_rd_data_2410;	// matmul/matmul-hw.mlir:15278:36, :15560:27, :15574:13
  assign c_i_k_9_i_j_2 = _T_3098;	// matmul/matmul-hw.mlir:15576:5
  //PROBE: c_i_k_9_i_j_2	// matmul/matmul-hw.mlir:15577:5
  assign _T_1166 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15578:13
  assign _T_1165 = _T_2874 ? _T_3098 : 32'bx;	// matmul/matmul-hw.mlir:9200:19, :15579:13
  localparam [3:0] _T_3100 = 4'h0;	// matmul/matmul-hw.mlir:15582:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15583:5
    if (rst)	// matmul/matmul-hw.mlir:15583:5
      i_k_next_3099 <= _T_3100;	// matmul/matmul-hw.mlir:15586:7
    else	// matmul/matmul-hw.mlir:15583:5
      i_k_next_3099 <= i_k_next_3096;	// matmul/matmul-hw.mlir:15551:13, :15584:7
  end // always @(posedge)
  assign _T_1164 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15588:13
  assign _T_1163 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15589:13
  mult mult_inst42 (	// matmul/matmul-hw.mlir:15590:27
    .a      (A_reg_bank42_p0_rd_data),	// matmul/matmul-hw.mlir:12257:32
    .b      (_T_2616),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst42_result)
  );
  assign _T_1162 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15591:13
  assign a_i_k_10_i_j_2 = A_reg_bank42_p0_rd_data;	// matmul/matmul-hw.mlir:12257:32, :15593:5
  //PROBE: a_i_k_10_i_j_2	// matmul/matmul-hw.mlir:15594:5
  assign b_i_k_10_i_j_2 = _T_2616;	// matmul/matmul-hw.mlir:15596:5
  //PROBE: b_i_k_10_i_j_2	// matmul/matmul-hw.mlir:15597:5
  assign c_prev_i_k_10_i_j_2 = C_reg_bank10_p0_rd_data_2409;	// matmul/matmul-hw.mlir:15279:37, :15599:5
  //PROBE: c_prev_i_k_10_i_j_2	// matmul/matmul-hw.mlir:15600:5
  assign tk_i_k_10_i_j_2 = _T_2841;	// matmul/matmul-hw.mlir:15602:5
  //PROBE: tk_i_k_10_i_j_2	// matmul/matmul-hw.mlir:15603:5
  wire [31:0] _T_3101 = mult_inst42_result + C_reg_bank10_p0_rd_data_2409;	// matmul/matmul-hw.mlir:15279:37, :15590:27, :15604:13
  assign c_i_k_10_i_j_2 = _T_3101;	// matmul/matmul-hw.mlir:15606:5
  //PROBE: c_i_k_10_i_j_2	// matmul/matmul-hw.mlir:15607:5
  assign _T_1161 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15608:13
  assign _T_1160 = _T_2885 ? _T_3101 : 32'bx;	// matmul/matmul-hw.mlir:9195:19, :15609:13
  localparam [3:0] _T_3103 = 4'h0;	// matmul/matmul-hw.mlir:15612:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15613:5
    if (rst)	// matmul/matmul-hw.mlir:15613:5
      i_k_next_3102 <= _T_3103;	// matmul/matmul-hw.mlir:15616:7
    else	// matmul/matmul-hw.mlir:15613:5
      i_k_next_3102 <= i_k_next_3099;	// matmul/matmul-hw.mlir:15581:13, :15614:7
  end // always @(posedge)
  assign _T_1159 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15618:13
  assign _T_1158 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15619:13
  mult mult_inst43 (	// matmul/matmul-hw.mlir:15620:27
    .a      (A_reg_bank43_p0_rd_data),	// matmul/matmul-hw.mlir:12258:32
    .b      (_T_2632),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst43_result)
  );
  assign _T_1157 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15621:13
  assign a_i_k_11_i_j_2 = A_reg_bank43_p0_rd_data;	// matmul/matmul-hw.mlir:12258:32, :15623:5
  //PROBE: a_i_k_11_i_j_2	// matmul/matmul-hw.mlir:15624:5
  assign b_i_k_11_i_j_2 = _T_2632;	// matmul/matmul-hw.mlir:15626:5
  //PROBE: b_i_k_11_i_j_2	// matmul/matmul-hw.mlir:15627:5
  assign c_prev_i_k_11_i_j_2 = C_reg_bank11_p0_rd_data_2408;	// matmul/matmul-hw.mlir:15280:37, :15629:5
  //PROBE: c_prev_i_k_11_i_j_2	// matmul/matmul-hw.mlir:15630:5
  assign tk_i_k_11_i_j_2 = _T_2852;	// matmul/matmul-hw.mlir:15632:5
  //PROBE: tk_i_k_11_i_j_2	// matmul/matmul-hw.mlir:15633:5
  wire [31:0] _T_3104 = mult_inst43_result + C_reg_bank11_p0_rd_data_2408;	// matmul/matmul-hw.mlir:15280:37, :15620:27, :15634:13
  assign c_i_k_11_i_j_2 = _T_3104;	// matmul/matmul-hw.mlir:15636:5
  //PROBE: c_i_k_11_i_j_2	// matmul/matmul-hw.mlir:15637:5
  assign _T_1156 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15638:13
  assign _T_1155 = _T_2892 ? _T_3104 : 32'bx;	// matmul/matmul-hw.mlir:9190:19, :15639:13
  localparam [3:0] _T_3106 = 4'h0;	// matmul/matmul-hw.mlir:15642:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15643:5
    if (rst)	// matmul/matmul-hw.mlir:15643:5
      i_k_next_3105 <= _T_3106;	// matmul/matmul-hw.mlir:15646:7
    else	// matmul/matmul-hw.mlir:15643:5
      i_k_next_3105 <= i_k_next_3102;	// matmul/matmul-hw.mlir:15611:13, :15644:7
  end // always @(posedge)
  assign _T_1154 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15648:13
  assign _T_1153 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15649:13
  mult mult_inst44 (	// matmul/matmul-hw.mlir:15650:27
    .a      (A_reg_bank44_p0_rd_data),	// matmul/matmul-hw.mlir:12259:32
    .b      (_T_2648),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst44_result)
  );
  assign _T_1152 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15651:13
  assign a_i_k_12_i_j_2 = A_reg_bank44_p0_rd_data;	// matmul/matmul-hw.mlir:12259:32, :15653:5
  //PROBE: a_i_k_12_i_j_2	// matmul/matmul-hw.mlir:15654:5
  assign b_i_k_12_i_j_2 = _T_2648;	// matmul/matmul-hw.mlir:15656:5
  //PROBE: b_i_k_12_i_j_2	// matmul/matmul-hw.mlir:15657:5
  assign c_prev_i_k_12_i_j_2 = C_reg_bank12_p0_rd_data_2407;	// matmul/matmul-hw.mlir:15281:37, :15659:5
  //PROBE: c_prev_i_k_12_i_j_2	// matmul/matmul-hw.mlir:15660:5
  assign tk_i_k_12_i_j_2 = _T_2863;	// matmul/matmul-hw.mlir:15662:5
  //PROBE: tk_i_k_12_i_j_2	// matmul/matmul-hw.mlir:15663:5
  wire [31:0] _T_3107 = mult_inst44_result + C_reg_bank12_p0_rd_data_2407;	// matmul/matmul-hw.mlir:15281:37, :15650:27, :15664:13
  assign c_i_k_12_i_j_2 = _T_3107;	// matmul/matmul-hw.mlir:15666:5
  //PROBE: c_i_k_12_i_j_2	// matmul/matmul-hw.mlir:15667:5
  assign _T_1151 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15668:13
  assign _T_1150 = _T_2897 ? _T_3107 : 32'bx;	// matmul/matmul-hw.mlir:9185:19, :15669:13
  localparam [3:0] _T_3109 = 4'h0;	// matmul/matmul-hw.mlir:15672:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15673:5
    if (rst)	// matmul/matmul-hw.mlir:15673:5
      i_k_next_3108 <= _T_3109;	// matmul/matmul-hw.mlir:15676:7
    else	// matmul/matmul-hw.mlir:15673:5
      i_k_next_3108 <= i_k_next_3105;	// matmul/matmul-hw.mlir:15641:13, :15674:7
  end // always @(posedge)
  assign _T_1149 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15678:13
  assign _T_1148 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15679:13
  mult mult_inst45 (	// matmul/matmul-hw.mlir:15680:27
    .a      (A_reg_bank45_p0_rd_data),	// matmul/matmul-hw.mlir:12260:32
    .b      (_T_2664),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst45_result)
  );
  assign _T_1147 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15681:13
  assign a_i_k_13_i_j_2 = A_reg_bank45_p0_rd_data;	// matmul/matmul-hw.mlir:12260:32, :15683:5
  //PROBE: a_i_k_13_i_j_2	// matmul/matmul-hw.mlir:15684:5
  assign b_i_k_13_i_j_2 = _T_2664;	// matmul/matmul-hw.mlir:15686:5
  //PROBE: b_i_k_13_i_j_2	// matmul/matmul-hw.mlir:15687:5
  assign c_prev_i_k_13_i_j_2 = C_reg_bank13_p0_rd_data_2406;	// matmul/matmul-hw.mlir:15282:37, :15689:5
  //PROBE: c_prev_i_k_13_i_j_2	// matmul/matmul-hw.mlir:15690:5
  assign tk_i_k_13_i_j_2 = _T_2874;	// matmul/matmul-hw.mlir:15692:5
  //PROBE: tk_i_k_13_i_j_2	// matmul/matmul-hw.mlir:15693:5
  wire [31:0] _T_3110 = mult_inst45_result + C_reg_bank13_p0_rd_data_2406;	// matmul/matmul-hw.mlir:15282:37, :15680:27, :15694:13
  assign c_i_k_13_i_j_2 = _T_3110;	// matmul/matmul-hw.mlir:15696:5
  //PROBE: c_i_k_13_i_j_2	// matmul/matmul-hw.mlir:15697:5
  assign _T_1146 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15698:13
  assign _T_1145 = _T_2902 ? _T_3110 : 32'bx;	// matmul/matmul-hw.mlir:9180:19, :15699:13
  localparam [3:0] _T_3112 = 4'h0;	// matmul/matmul-hw.mlir:15702:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15703:5
    if (rst)	// matmul/matmul-hw.mlir:15703:5
      i_k_next_3111 <= _T_3112;	// matmul/matmul-hw.mlir:15706:7
    else	// matmul/matmul-hw.mlir:15703:5
      i_k_next_3111 <= i_k_next_3108;	// matmul/matmul-hw.mlir:15671:13, :15704:7
  end // always @(posedge)
  assign _T_1144 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15708:13
  assign _T_1143 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15709:13
  mult mult_inst46 (	// matmul/matmul-hw.mlir:15710:27
    .a      (A_reg_bank46_p0_rd_data),	// matmul/matmul-hw.mlir:12261:32
    .b      (_T_2680),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst46_result)
  );
  assign _T_1142 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15711:13
  assign a_i_k_14_i_j_2 = A_reg_bank46_p0_rd_data;	// matmul/matmul-hw.mlir:12261:32, :15713:5
  //PROBE: a_i_k_14_i_j_2	// matmul/matmul-hw.mlir:15714:5
  assign b_i_k_14_i_j_2 = _T_2680;	// matmul/matmul-hw.mlir:15716:5
  //PROBE: b_i_k_14_i_j_2	// matmul/matmul-hw.mlir:15717:5
  assign c_prev_i_k_14_i_j_2 = C_reg_bank14_p0_rd_data_2405;	// matmul/matmul-hw.mlir:15283:37, :15719:5
  //PROBE: c_prev_i_k_14_i_j_2	// matmul/matmul-hw.mlir:15720:5
  assign tk_i_k_14_i_j_2 = _T_2885;	// matmul/matmul-hw.mlir:15722:5
  //PROBE: tk_i_k_14_i_j_2	// matmul/matmul-hw.mlir:15723:5
  wire [31:0] _T_3113 = mult_inst46_result + C_reg_bank14_p0_rd_data_2405;	// matmul/matmul-hw.mlir:15283:37, :15710:27, :15724:13
  assign c_i_k_14_i_j_2 = _T_3113;	// matmul/matmul-hw.mlir:15726:5
  //PROBE: c_i_k_14_i_j_2	// matmul/matmul-hw.mlir:15727:5
  assign _T_1141 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15728:13
  assign _T_1140 = _T_2907 ? _T_3113 : 32'bx;	// matmul/matmul-hw.mlir:9175:19, :15729:13
  localparam [3:0] _T_3115 = 4'h0;	// matmul/matmul-hw.mlir:15732:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15733:5
    if (rst)	// matmul/matmul-hw.mlir:15733:5
      i_k_next_3114 <= _T_3115;	// matmul/matmul-hw.mlir:15736:7
    else	// matmul/matmul-hw.mlir:15733:5
      i_k_next_3114 <= i_k_next_3111;	// matmul/matmul-hw.mlir:15701:13, :15734:7
  end // always @(posedge)
  assign _T_1139 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15738:13
  assign _T_1138 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15739:13
  mult mult_inst47 (	// matmul/matmul-hw.mlir:15740:27
    .a      (A_reg_bank47_p0_rd_data),	// matmul/matmul-hw.mlir:12262:32
    .b      (_T_2696),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst47_result)
  );
  assign _T_1137 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15741:13
  assign a_i_k_15_i_j_2 = A_reg_bank47_p0_rd_data;	// matmul/matmul-hw.mlir:12262:32, :15743:5
  //PROBE: a_i_k_15_i_j_2	// matmul/matmul-hw.mlir:15744:5
  assign b_i_k_15_i_j_2 = _T_2696;	// matmul/matmul-hw.mlir:15746:5
  //PROBE: b_i_k_15_i_j_2	// matmul/matmul-hw.mlir:15747:5
  assign c_prev_i_k_15_i_j_2 = C_reg_bank15_p0_rd_data_2404;	// matmul/matmul-hw.mlir:15284:37, :15749:5
  //PROBE: c_prev_i_k_15_i_j_2	// matmul/matmul-hw.mlir:15750:5
  assign tk_i_k_15_i_j_2 = _T_2892;	// matmul/matmul-hw.mlir:15752:5
  //PROBE: tk_i_k_15_i_j_2	// matmul/matmul-hw.mlir:15753:5
  wire [31:0] _T_3116 = mult_inst47_result + C_reg_bank15_p0_rd_data_2404;	// matmul/matmul-hw.mlir:15284:37, :15740:27, :15754:13
  assign c_i_k_15_i_j_2 = _T_3116;	// matmul/matmul-hw.mlir:15756:5
  //PROBE: c_i_k_15_i_j_2	// matmul/matmul-hw.mlir:15757:5
  assign _T_1136 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15758:13
  assign _T_1135 = _T_2912 ? _T_3116 : 32'bx;	// matmul/matmul-hw.mlir:9170:19, :15759:13
  localparam [3:0] _T_3118 = 4'h0;	// matmul/matmul-hw.mlir:15762:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15763:5
    if (rst)	// matmul/matmul-hw.mlir:15763:5
      i_k_next_3117 <= _T_3118;	// matmul/matmul-hw.mlir:15766:7
    else	// matmul/matmul-hw.mlir:15763:5
      i_k_next_3117 <= i_k_next_3114;	// matmul/matmul-hw.mlir:15731:13, :15764:7
  end // always @(posedge)
  assign _T_1134 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15768:13
  wire [3:0][3:0] _T_3120 = i_delayed_3119;	// matmul/matmul-hw.mlir:15770:13
  wire [3:0][3:0] _T_3121 = {_T_3120[2'h0+:3], {{i_k_next_3117}}};	// matmul/matmul-hw.mlir:15761:13, :15771:19, :15772:13, :15773:13, :15774:13
  wire [3:0][3:0] _T_3122 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:15775:19, :15776:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15777:5
    if (rst)	// matmul/matmul-hw.mlir:15777:5
      i_delayed_3119 <= _T_3122;	// matmul/matmul-hw.mlir:15780:7
    else	// matmul/matmul-hw.mlir:15777:5
      i_delayed_3119 <= _T_3121;	// matmul/matmul-hw.mlir:15778:7
  end // always @(posedge)
  assign _T_1133 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15784:13
  assign _T_1132 = _T_2917 ? i_delayed_3119[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:9167:18, :15770:13, :15782:20, :15783:13, :15785:13
  assign _T_1131 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15786:13
  assign _T_1130 = _T_2917 ? C_reg_bank16_p0_rd_data_2403 : 32'bx;	// matmul/matmul-hw.mlir:9165:19, :15285:37, :15787:13
  localparam [3:0] _T_3124 = 4'h0;	// matmul/matmul-hw.mlir:15790:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15791:5
    if (rst)	// matmul/matmul-hw.mlir:15791:5
      i_j_next_3123 <= _T_3124;	// matmul/matmul-hw.mlir:15794:7
    else	// matmul/matmul-hw.mlir:15791:5
      i_j_next_3123 <= i_j_next_3052;	// matmul/matmul-hw.mlir:15194:13, :15792:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3125 (	// matmul/matmul-hw.mlir:15864:36
    .p0_rd_en   (_T_1125),	// matmul/matmul-hw.mlir:15886:13
    .p1_wr_en   (_T_1129),	// matmul/matmul-hw.mlir:15881:13
    .p1_wr_data (_T_1128),	// matmul/matmul-hw.mlir:15882:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2402)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3126 (	// matmul/matmul-hw.mlir:15865:36
    .p0_rd_en   (_T_1120),	// matmul/matmul-hw.mlir:15916:13
    .p1_wr_en   (_T_1124),	// matmul/matmul-hw.mlir:15903:13
    .p1_wr_data (_T_1123),	// matmul/matmul-hw.mlir:15904:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2401)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3127 (	// matmul/matmul-hw.mlir:15866:36
    .p0_rd_en   (_T_1115),	// matmul/matmul-hw.mlir:15946:13
    .p1_wr_en   (_T_1119),	// matmul/matmul-hw.mlir:15933:13
    .p1_wr_data (_T_1118),	// matmul/matmul-hw.mlir:15934:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2400)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3128 (	// matmul/matmul-hw.mlir:15867:36
    .p0_rd_en   (_T_1110),	// matmul/matmul-hw.mlir:15976:13
    .p1_wr_en   (_T_1114),	// matmul/matmul-hw.mlir:15963:13
    .p1_wr_data (_T_1113),	// matmul/matmul-hw.mlir:15964:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2399)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3129 (	// matmul/matmul-hw.mlir:15868:36
    .p0_rd_en   (_T_1105),	// matmul/matmul-hw.mlir:16006:13
    .p1_wr_en   (_T_1109),	// matmul/matmul-hw.mlir:15993:13
    .p1_wr_data (_T_1108),	// matmul/matmul-hw.mlir:15994:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2398)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3130 (	// matmul/matmul-hw.mlir:15869:36
    .p0_rd_en   (_T_1100),	// matmul/matmul-hw.mlir:16036:13
    .p1_wr_en   (_T_1104),	// matmul/matmul-hw.mlir:16023:13
    .p1_wr_data (_T_1103),	// matmul/matmul-hw.mlir:16024:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2397)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3131 (	// matmul/matmul-hw.mlir:15870:36
    .p0_rd_en   (_T_1095),	// matmul/matmul-hw.mlir:16066:13
    .p1_wr_en   (_T_1099),	// matmul/matmul-hw.mlir:16053:13
    .p1_wr_data (_T_1098),	// matmul/matmul-hw.mlir:16054:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2396)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3132 (	// matmul/matmul-hw.mlir:15871:36
    .p0_rd_en   (_T_1090),	// matmul/matmul-hw.mlir:16096:13
    .p1_wr_en   (_T_1094),	// matmul/matmul-hw.mlir:16083:13
    .p1_wr_data (_T_1093),	// matmul/matmul-hw.mlir:16084:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2395)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3133 (	// matmul/matmul-hw.mlir:15872:36
    .p0_rd_en   (_T_1085),	// matmul/matmul-hw.mlir:16126:13
    .p1_wr_en   (_T_1089),	// matmul/matmul-hw.mlir:16113:13
    .p1_wr_data (_T_1088),	// matmul/matmul-hw.mlir:16114:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2394)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3134 (	// matmul/matmul-hw.mlir:15873:36
    .p0_rd_en   (_T_1080),	// matmul/matmul-hw.mlir:16156:13
    .p1_wr_en   (_T_1084),	// matmul/matmul-hw.mlir:16143:13
    .p1_wr_data (_T_1083),	// matmul/matmul-hw.mlir:16144:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2393)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3135 (	// matmul/matmul-hw.mlir:15874:37
    .p0_rd_en   (_T_1075),	// matmul/matmul-hw.mlir:16186:13
    .p1_wr_en   (_T_1079),	// matmul/matmul-hw.mlir:16173:13
    .p1_wr_data (_T_1078),	// matmul/matmul-hw.mlir:16174:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2392)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3136 (	// matmul/matmul-hw.mlir:15875:37
    .p0_rd_en   (_T_1070),	// matmul/matmul-hw.mlir:16216:13
    .p1_wr_en   (_T_1074),	// matmul/matmul-hw.mlir:16203:13
    .p1_wr_data (_T_1073),	// matmul/matmul-hw.mlir:16204:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2391)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3137 (	// matmul/matmul-hw.mlir:15876:37
    .p0_rd_en   (_T_1065),	// matmul/matmul-hw.mlir:16246:13
    .p1_wr_en   (_T_1069),	// matmul/matmul-hw.mlir:16233:13
    .p1_wr_data (_T_1068),	// matmul/matmul-hw.mlir:16234:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2390)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3138 (	// matmul/matmul-hw.mlir:15877:37
    .p0_rd_en   (_T_1060),	// matmul/matmul-hw.mlir:16276:13
    .p1_wr_en   (_T_1064),	// matmul/matmul-hw.mlir:16263:13
    .p1_wr_data (_T_1063),	// matmul/matmul-hw.mlir:16264:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2389)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3139 (	// matmul/matmul-hw.mlir:15878:37
    .p0_rd_en   (_T_1055),	// matmul/matmul-hw.mlir:16306:13
    .p1_wr_en   (_T_1059),	// matmul/matmul-hw.mlir:16293:13
    .p1_wr_data (_T_1058),	// matmul/matmul-hw.mlir:16294:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2388)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3140 (	// matmul/matmul-hw.mlir:15879:37
    .p0_rd_en   (_T_1050),	// matmul/matmul-hw.mlir:16336:13
    .p1_wr_en   (_T_1054),	// matmul/matmul-hw.mlir:16323:13
    .p1_wr_data (_T_1053),	// matmul/matmul-hw.mlir:16324:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2387)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3141 (	// matmul/matmul-hw.mlir:15880:37
    .p0_rd_en   (_T_1047),	// matmul/matmul-hw.mlir:16363:13
    .p1_wr_en   (_T_1049),	// matmul/matmul-hw.mlir:16353:13
    .p1_wr_data (_T_1048),	// matmul/matmul-hw.mlir:16354:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2386)
  );
  assign _T_1129 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15881:13
  assign _T_1128 = _T_2775 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :9163:19, :15882:13
  assign _T_1127 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15883:13
  assign _T_1126 = _T_2764 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15884:13
  mult mult_inst48 (	// matmul/matmul-hw.mlir:15885:27
    .a      (A_reg_bank48_p0_rd_data),	// matmul/matmul-hw.mlir:12263:32
    .b      (_T_2457),
    .t      (_T_2764),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst48_result)
  );
  assign _T_1125 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15886:13
  assign a_i_k_0_i_j_3 = A_reg_bank48_p0_rd_data;	// matmul/matmul-hw.mlir:12263:32, :15888:5
  //PROBE: a_i_k_0_i_j_3	// matmul/matmul-hw.mlir:15889:5
  assign b_i_k_0_i_j_3 = _T_2457;	// matmul/matmul-hw.mlir:15891:5
  //PROBE: b_i_k_0_i_j_3	// matmul/matmul-hw.mlir:15892:5
  assign c_prev_i_k_0_i_j_3 = C_reg_bank0_p0_rd_data_2402;	// matmul/matmul-hw.mlir:15864:36, :15894:5
  //PROBE: c_prev_i_k_0_i_j_3	// matmul/matmul-hw.mlir:15895:5
  assign tk_i_k_0_i_j_3 = _T_2742;	// matmul/matmul-hw.mlir:15897:5
  //PROBE: tk_i_k_0_i_j_3	// matmul/matmul-hw.mlir:15898:5
  wire [31:0] _T_3142 = mult_inst48_result + C_reg_bank0_p0_rd_data_2402;	// matmul/matmul-hw.mlir:15864:36, :15885:27, :15899:13
  assign c_i_k_0_i_j_3 = _T_3142;	// matmul/matmul-hw.mlir:15901:5
  //PROBE: c_i_k_0_i_j_3	// matmul/matmul-hw.mlir:15902:5
  assign _T_1124 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15903:13
  assign _T_1123 = _T_2786 ? _T_3142 : 32'bx;	// matmul/matmul-hw.mlir:9158:19, :15904:13
  localparam [3:0] _T_3144 = 4'h0;	// matmul/matmul-hw.mlir:15907:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15908:5
    if (rst)	// matmul/matmul-hw.mlir:15908:5
      i_k_next_3143 <= _T_3144;	// matmul/matmul-hw.mlir:15911:7
    else	// matmul/matmul-hw.mlir:15908:5
      i_k_next_3143 <= i_j_next_3123;	// matmul/matmul-hw.mlir:15789:13, :15909:7
  end // always @(posedge)
  assign _T_1122 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15913:13
  assign _T_1121 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15914:13
  mult mult_inst49 (	// matmul/matmul-hw.mlir:15915:27
    .a      (A_reg_bank49_p0_rd_data),	// matmul/matmul-hw.mlir:12264:32
    .b      (_T_2473),
    .t      (_T_2775),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst49_result)
  );
  assign _T_1120 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15916:13
  assign a_i_k_1_i_j_3 = A_reg_bank49_p0_rd_data;	// matmul/matmul-hw.mlir:12264:32, :15918:5
  //PROBE: a_i_k_1_i_j_3	// matmul/matmul-hw.mlir:15919:5
  assign b_i_k_1_i_j_3 = _T_2473;	// matmul/matmul-hw.mlir:15921:5
  //PROBE: b_i_k_1_i_j_3	// matmul/matmul-hw.mlir:15922:5
  assign c_prev_i_k_1_i_j_3 = C_reg_bank1_p0_rd_data_2401;	// matmul/matmul-hw.mlir:15865:36, :15924:5
  //PROBE: c_prev_i_k_1_i_j_3	// matmul/matmul-hw.mlir:15925:5
  assign tk_i_k_1_i_j_3 = _T_2753;	// matmul/matmul-hw.mlir:15927:5
  //PROBE: tk_i_k_1_i_j_3	// matmul/matmul-hw.mlir:15928:5
  wire [31:0] _T_3145 = mult_inst49_result + C_reg_bank1_p0_rd_data_2401;	// matmul/matmul-hw.mlir:15865:36, :15915:27, :15929:13
  assign c_i_k_1_i_j_3 = _T_3145;	// matmul/matmul-hw.mlir:15931:5
  //PROBE: c_i_k_1_i_j_3	// matmul/matmul-hw.mlir:15932:5
  assign _T_1119 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15933:13
  assign _T_1118 = _T_2797 ? _T_3145 : 32'bx;	// matmul/matmul-hw.mlir:9153:19, :15934:13
  localparam [3:0] _T_3147 = 4'h0;	// matmul/matmul-hw.mlir:15937:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15938:5
    if (rst)	// matmul/matmul-hw.mlir:15938:5
      i_k_next_3146 <= _T_3147;	// matmul/matmul-hw.mlir:15941:7
    else	// matmul/matmul-hw.mlir:15938:5
      i_k_next_3146 <= i_k_next_3143;	// matmul/matmul-hw.mlir:15906:13, :15939:7
  end // always @(posedge)
  assign _T_1117 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15943:13
  assign _T_1116 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15944:13
  mult mult_inst50 (	// matmul/matmul-hw.mlir:15945:27
    .a      (A_reg_bank50_p0_rd_data),	// matmul/matmul-hw.mlir:12265:32
    .b      (_T_2489),
    .t      (_T_2786),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst50_result)
  );
  assign _T_1115 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15946:13
  assign a_i_k_2_i_j_3 = A_reg_bank50_p0_rd_data;	// matmul/matmul-hw.mlir:12265:32, :15948:5
  //PROBE: a_i_k_2_i_j_3	// matmul/matmul-hw.mlir:15949:5
  assign b_i_k_2_i_j_3 = _T_2489;	// matmul/matmul-hw.mlir:15951:5
  //PROBE: b_i_k_2_i_j_3	// matmul/matmul-hw.mlir:15952:5
  assign c_prev_i_k_2_i_j_3 = C_reg_bank2_p0_rd_data_2400;	// matmul/matmul-hw.mlir:15866:36, :15954:5
  //PROBE: c_prev_i_k_2_i_j_3	// matmul/matmul-hw.mlir:15955:5
  assign tk_i_k_2_i_j_3 = _T_2764;	// matmul/matmul-hw.mlir:15957:5
  //PROBE: tk_i_k_2_i_j_3	// matmul/matmul-hw.mlir:15958:5
  wire [31:0] _T_3148 = mult_inst50_result + C_reg_bank2_p0_rd_data_2400;	// matmul/matmul-hw.mlir:15866:36, :15945:27, :15959:13
  assign c_i_k_2_i_j_3 = _T_3148;	// matmul/matmul-hw.mlir:15961:5
  //PROBE: c_i_k_2_i_j_3	// matmul/matmul-hw.mlir:15962:5
  assign _T_1114 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15963:13
  assign _T_1113 = _T_2808 ? _T_3148 : 32'bx;	// matmul/matmul-hw.mlir:9148:19, :15964:13
  localparam [3:0] _T_3150 = 4'h0;	// matmul/matmul-hw.mlir:15967:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15968:5
    if (rst)	// matmul/matmul-hw.mlir:15968:5
      i_k_next_3149 <= _T_3150;	// matmul/matmul-hw.mlir:15971:7
    else	// matmul/matmul-hw.mlir:15968:5
      i_k_next_3149 <= i_k_next_3146;	// matmul/matmul-hw.mlir:15936:13, :15969:7
  end // always @(posedge)
  assign _T_1112 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15973:13
  assign _T_1111 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15974:13
  mult mult_inst51 (	// matmul/matmul-hw.mlir:15975:27
    .a      (A_reg_bank51_p0_rd_data),	// matmul/matmul-hw.mlir:12266:32
    .b      (_T_2505),
    .t      (_T_2797),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst51_result)
  );
  assign _T_1110 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15976:13
  assign a_i_k_3_i_j_3 = A_reg_bank51_p0_rd_data;	// matmul/matmul-hw.mlir:12266:32, :15978:5
  //PROBE: a_i_k_3_i_j_3	// matmul/matmul-hw.mlir:15979:5
  assign b_i_k_3_i_j_3 = _T_2505;	// matmul/matmul-hw.mlir:15981:5
  //PROBE: b_i_k_3_i_j_3	// matmul/matmul-hw.mlir:15982:5
  assign c_prev_i_k_3_i_j_3 = C_reg_bank3_p0_rd_data_2399;	// matmul/matmul-hw.mlir:15867:36, :15984:5
  //PROBE: c_prev_i_k_3_i_j_3	// matmul/matmul-hw.mlir:15985:5
  assign tk_i_k_3_i_j_3 = _T_2775;	// matmul/matmul-hw.mlir:15987:5
  //PROBE: tk_i_k_3_i_j_3	// matmul/matmul-hw.mlir:15988:5
  wire [31:0] _T_3151 = mult_inst51_result + C_reg_bank3_p0_rd_data_2399;	// matmul/matmul-hw.mlir:15867:36, :15975:27, :15989:13
  assign c_i_k_3_i_j_3 = _T_3151;	// matmul/matmul-hw.mlir:15991:5
  //PROBE: c_i_k_3_i_j_3	// matmul/matmul-hw.mlir:15992:5
  assign _T_1109 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :15993:13
  assign _T_1108 = _T_2819 ? _T_3151 : 32'bx;	// matmul/matmul-hw.mlir:9143:19, :15994:13
  localparam [3:0] _T_3153 = 4'h0;	// matmul/matmul-hw.mlir:15997:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:15998:5
    if (rst)	// matmul/matmul-hw.mlir:15998:5
      i_k_next_3152 <= _T_3153;	// matmul/matmul-hw.mlir:16001:7
    else	// matmul/matmul-hw.mlir:15998:5
      i_k_next_3152 <= i_k_next_3149;	// matmul/matmul-hw.mlir:15966:13, :15999:7
  end // always @(posedge)
  assign _T_1107 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16003:13
  assign _T_1106 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16004:13
  mult mult_inst52 (	// matmul/matmul-hw.mlir:16005:27
    .a      (A_reg_bank52_p0_rd_data),	// matmul/matmul-hw.mlir:12267:32
    .b      (_T_2521),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst52_result)
  );
  assign _T_1105 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16006:13
  assign a_i_k_4_i_j_3 = A_reg_bank52_p0_rd_data;	// matmul/matmul-hw.mlir:12267:32, :16008:5
  //PROBE: a_i_k_4_i_j_3	// matmul/matmul-hw.mlir:16009:5
  assign b_i_k_4_i_j_3 = _T_2521;	// matmul/matmul-hw.mlir:16011:5
  //PROBE: b_i_k_4_i_j_3	// matmul/matmul-hw.mlir:16012:5
  assign c_prev_i_k_4_i_j_3 = C_reg_bank4_p0_rd_data_2398;	// matmul/matmul-hw.mlir:15868:36, :16014:5
  //PROBE: c_prev_i_k_4_i_j_3	// matmul/matmul-hw.mlir:16015:5
  assign tk_i_k_4_i_j_3 = _T_2786;	// matmul/matmul-hw.mlir:16017:5
  //PROBE: tk_i_k_4_i_j_3	// matmul/matmul-hw.mlir:16018:5
  wire [31:0] _T_3154 = mult_inst52_result + C_reg_bank4_p0_rd_data_2398;	// matmul/matmul-hw.mlir:15868:36, :16005:27, :16019:13
  assign c_i_k_4_i_j_3 = _T_3154;	// matmul/matmul-hw.mlir:16021:5
  //PROBE: c_i_k_4_i_j_3	// matmul/matmul-hw.mlir:16022:5
  assign _T_1104 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16023:13
  assign _T_1103 = _T_2830 ? _T_3154 : 32'bx;	// matmul/matmul-hw.mlir:9138:19, :16024:13
  localparam [3:0] _T_3156 = 4'h0;	// matmul/matmul-hw.mlir:16027:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16028:5
    if (rst)	// matmul/matmul-hw.mlir:16028:5
      i_k_next_3155 <= _T_3156;	// matmul/matmul-hw.mlir:16031:7
    else	// matmul/matmul-hw.mlir:16028:5
      i_k_next_3155 <= i_k_next_3152;	// matmul/matmul-hw.mlir:15996:13, :16029:7
  end // always @(posedge)
  assign _T_1102 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16033:13
  assign _T_1101 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16034:13
  mult mult_inst53 (	// matmul/matmul-hw.mlir:16035:27
    .a      (A_reg_bank53_p0_rd_data),	// matmul/matmul-hw.mlir:12268:32
    .b      (_T_2537),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst53_result)
  );
  assign _T_1100 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16036:13
  assign a_i_k_5_i_j_3 = A_reg_bank53_p0_rd_data;	// matmul/matmul-hw.mlir:12268:32, :16038:5
  //PROBE: a_i_k_5_i_j_3	// matmul/matmul-hw.mlir:16039:5
  assign b_i_k_5_i_j_3 = _T_2537;	// matmul/matmul-hw.mlir:16041:5
  //PROBE: b_i_k_5_i_j_3	// matmul/matmul-hw.mlir:16042:5
  assign c_prev_i_k_5_i_j_3 = C_reg_bank5_p0_rd_data_2397;	// matmul/matmul-hw.mlir:15869:36, :16044:5
  //PROBE: c_prev_i_k_5_i_j_3	// matmul/matmul-hw.mlir:16045:5
  assign tk_i_k_5_i_j_3 = _T_2797;	// matmul/matmul-hw.mlir:16047:5
  //PROBE: tk_i_k_5_i_j_3	// matmul/matmul-hw.mlir:16048:5
  wire [31:0] _T_3157 = mult_inst53_result + C_reg_bank5_p0_rd_data_2397;	// matmul/matmul-hw.mlir:15869:36, :16035:27, :16049:13
  assign c_i_k_5_i_j_3 = _T_3157;	// matmul/matmul-hw.mlir:16051:5
  //PROBE: c_i_k_5_i_j_3	// matmul/matmul-hw.mlir:16052:5
  assign _T_1099 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16053:13
  assign _T_1098 = _T_2841 ? _T_3157 : 32'bx;	// matmul/matmul-hw.mlir:9133:19, :16054:13
  localparam [3:0] _T_3159 = 4'h0;	// matmul/matmul-hw.mlir:16057:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16058:5
    if (rst)	// matmul/matmul-hw.mlir:16058:5
      i_k_next_3158 <= _T_3159;	// matmul/matmul-hw.mlir:16061:7
    else	// matmul/matmul-hw.mlir:16058:5
      i_k_next_3158 <= i_k_next_3155;	// matmul/matmul-hw.mlir:16026:13, :16059:7
  end // always @(posedge)
  assign _T_1097 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16063:13
  assign _T_1096 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16064:13
  mult mult_inst54 (	// matmul/matmul-hw.mlir:16065:27
    .a      (A_reg_bank54_p0_rd_data),	// matmul/matmul-hw.mlir:12269:32
    .b      (_T_2553),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst54_result)
  );
  assign _T_1095 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16066:13
  assign a_i_k_6_i_j_3 = A_reg_bank54_p0_rd_data;	// matmul/matmul-hw.mlir:12269:32, :16068:5
  //PROBE: a_i_k_6_i_j_3	// matmul/matmul-hw.mlir:16069:5
  assign b_i_k_6_i_j_3 = _T_2553;	// matmul/matmul-hw.mlir:16071:5
  //PROBE: b_i_k_6_i_j_3	// matmul/matmul-hw.mlir:16072:5
  assign c_prev_i_k_6_i_j_3 = C_reg_bank6_p0_rd_data_2396;	// matmul/matmul-hw.mlir:15870:36, :16074:5
  //PROBE: c_prev_i_k_6_i_j_3	// matmul/matmul-hw.mlir:16075:5
  assign tk_i_k_6_i_j_3 = _T_2808;	// matmul/matmul-hw.mlir:16077:5
  //PROBE: tk_i_k_6_i_j_3	// matmul/matmul-hw.mlir:16078:5
  wire [31:0] _T_3160 = mult_inst54_result + C_reg_bank6_p0_rd_data_2396;	// matmul/matmul-hw.mlir:15870:36, :16065:27, :16079:13
  assign c_i_k_6_i_j_3 = _T_3160;	// matmul/matmul-hw.mlir:16081:5
  //PROBE: c_i_k_6_i_j_3	// matmul/matmul-hw.mlir:16082:5
  assign _T_1094 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16083:13
  assign _T_1093 = _T_2852 ? _T_3160 : 32'bx;	// matmul/matmul-hw.mlir:9128:19, :16084:13
  localparam [3:0] _T_3162 = 4'h0;	// matmul/matmul-hw.mlir:16087:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16088:5
    if (rst)	// matmul/matmul-hw.mlir:16088:5
      i_k_next_3161 <= _T_3162;	// matmul/matmul-hw.mlir:16091:7
    else	// matmul/matmul-hw.mlir:16088:5
      i_k_next_3161 <= i_k_next_3158;	// matmul/matmul-hw.mlir:16056:13, :16089:7
  end // always @(posedge)
  assign _T_1092 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16093:13
  assign _T_1091 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16094:13
  mult mult_inst55 (	// matmul/matmul-hw.mlir:16095:27
    .a      (A_reg_bank55_p0_rd_data),	// matmul/matmul-hw.mlir:12270:32
    .b      (_T_2569),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst55_result)
  );
  assign _T_1090 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16096:13
  assign a_i_k_7_i_j_3 = A_reg_bank55_p0_rd_data;	// matmul/matmul-hw.mlir:12270:32, :16098:5
  //PROBE: a_i_k_7_i_j_3	// matmul/matmul-hw.mlir:16099:5
  assign b_i_k_7_i_j_3 = _T_2569;	// matmul/matmul-hw.mlir:16101:5
  //PROBE: b_i_k_7_i_j_3	// matmul/matmul-hw.mlir:16102:5
  assign c_prev_i_k_7_i_j_3 = C_reg_bank7_p0_rd_data_2395;	// matmul/matmul-hw.mlir:15871:36, :16104:5
  //PROBE: c_prev_i_k_7_i_j_3	// matmul/matmul-hw.mlir:16105:5
  assign tk_i_k_7_i_j_3 = _T_2819;	// matmul/matmul-hw.mlir:16107:5
  //PROBE: tk_i_k_7_i_j_3	// matmul/matmul-hw.mlir:16108:5
  wire [31:0] _T_3163 = mult_inst55_result + C_reg_bank7_p0_rd_data_2395;	// matmul/matmul-hw.mlir:15871:36, :16095:27, :16109:13
  assign c_i_k_7_i_j_3 = _T_3163;	// matmul/matmul-hw.mlir:16111:5
  //PROBE: c_i_k_7_i_j_3	// matmul/matmul-hw.mlir:16112:5
  assign _T_1089 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16113:13
  assign _T_1088 = _T_2863 ? _T_3163 : 32'bx;	// matmul/matmul-hw.mlir:9123:19, :16114:13
  localparam [3:0] _T_3165 = 4'h0;	// matmul/matmul-hw.mlir:16117:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16118:5
    if (rst)	// matmul/matmul-hw.mlir:16118:5
      i_k_next_3164 <= _T_3165;	// matmul/matmul-hw.mlir:16121:7
    else	// matmul/matmul-hw.mlir:16118:5
      i_k_next_3164 <= i_k_next_3161;	// matmul/matmul-hw.mlir:16086:13, :16119:7
  end // always @(posedge)
  assign _T_1087 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16123:13
  assign _T_1086 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16124:13
  mult mult_inst56 (	// matmul/matmul-hw.mlir:16125:27
    .a      (A_reg_bank56_p0_rd_data),	// matmul/matmul-hw.mlir:12271:32
    .b      (_T_2585),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst56_result)
  );
  assign _T_1085 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16126:13
  assign a_i_k_8_i_j_3 = A_reg_bank56_p0_rd_data;	// matmul/matmul-hw.mlir:12271:32, :16128:5
  //PROBE: a_i_k_8_i_j_3	// matmul/matmul-hw.mlir:16129:5
  assign b_i_k_8_i_j_3 = _T_2585;	// matmul/matmul-hw.mlir:16131:5
  //PROBE: b_i_k_8_i_j_3	// matmul/matmul-hw.mlir:16132:5
  assign c_prev_i_k_8_i_j_3 = C_reg_bank8_p0_rd_data_2394;	// matmul/matmul-hw.mlir:15872:36, :16134:5
  //PROBE: c_prev_i_k_8_i_j_3	// matmul/matmul-hw.mlir:16135:5
  assign tk_i_k_8_i_j_3 = _T_2830;	// matmul/matmul-hw.mlir:16137:5
  //PROBE: tk_i_k_8_i_j_3	// matmul/matmul-hw.mlir:16138:5
  wire [31:0] _T_3166 = mult_inst56_result + C_reg_bank8_p0_rd_data_2394;	// matmul/matmul-hw.mlir:15872:36, :16125:27, :16139:13
  assign c_i_k_8_i_j_3 = _T_3166;	// matmul/matmul-hw.mlir:16141:5
  //PROBE: c_i_k_8_i_j_3	// matmul/matmul-hw.mlir:16142:5
  assign _T_1084 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16143:13
  assign _T_1083 = _T_2874 ? _T_3166 : 32'bx;	// matmul/matmul-hw.mlir:9118:19, :16144:13
  localparam [3:0] _T_3168 = 4'h0;	// matmul/matmul-hw.mlir:16147:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16148:5
    if (rst)	// matmul/matmul-hw.mlir:16148:5
      i_k_next_3167 <= _T_3168;	// matmul/matmul-hw.mlir:16151:7
    else	// matmul/matmul-hw.mlir:16148:5
      i_k_next_3167 <= i_k_next_3164;	// matmul/matmul-hw.mlir:16116:13, :16149:7
  end // always @(posedge)
  assign _T_1082 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16153:13
  assign _T_1081 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16154:13
  mult mult_inst57 (	// matmul/matmul-hw.mlir:16155:27
    .a      (A_reg_bank57_p0_rd_data),	// matmul/matmul-hw.mlir:12272:32
    .b      (_T_2601),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst57_result)
  );
  assign _T_1080 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16156:13
  assign a_i_k_9_i_j_3 = A_reg_bank57_p0_rd_data;	// matmul/matmul-hw.mlir:12272:32, :16158:5
  //PROBE: a_i_k_9_i_j_3	// matmul/matmul-hw.mlir:16159:5
  assign b_i_k_9_i_j_3 = _T_2601;	// matmul/matmul-hw.mlir:16161:5
  //PROBE: b_i_k_9_i_j_3	// matmul/matmul-hw.mlir:16162:5
  assign c_prev_i_k_9_i_j_3 = C_reg_bank9_p0_rd_data_2393;	// matmul/matmul-hw.mlir:15873:36, :16164:5
  //PROBE: c_prev_i_k_9_i_j_3	// matmul/matmul-hw.mlir:16165:5
  assign tk_i_k_9_i_j_3 = _T_2841;	// matmul/matmul-hw.mlir:16167:5
  //PROBE: tk_i_k_9_i_j_3	// matmul/matmul-hw.mlir:16168:5
  wire [31:0] _T_3169 = mult_inst57_result + C_reg_bank9_p0_rd_data_2393;	// matmul/matmul-hw.mlir:15873:36, :16155:27, :16169:13
  assign c_i_k_9_i_j_3 = _T_3169;	// matmul/matmul-hw.mlir:16171:5
  //PROBE: c_i_k_9_i_j_3	// matmul/matmul-hw.mlir:16172:5
  assign _T_1079 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16173:13
  assign _T_1078 = _T_2885 ? _T_3169 : 32'bx;	// matmul/matmul-hw.mlir:9113:19, :16174:13
  localparam [3:0] _T_3171 = 4'h0;	// matmul/matmul-hw.mlir:16177:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16178:5
    if (rst)	// matmul/matmul-hw.mlir:16178:5
      i_k_next_3170 <= _T_3171;	// matmul/matmul-hw.mlir:16181:7
    else	// matmul/matmul-hw.mlir:16178:5
      i_k_next_3170 <= i_k_next_3167;	// matmul/matmul-hw.mlir:16146:13, :16179:7
  end // always @(posedge)
  assign _T_1077 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16183:13
  assign _T_1076 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16184:13
  mult mult_inst58 (	// matmul/matmul-hw.mlir:16185:27
    .a      (A_reg_bank58_p0_rd_data),	// matmul/matmul-hw.mlir:12273:32
    .b      (_T_2617),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst58_result)
  );
  assign _T_1075 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16186:13
  assign a_i_k_10_i_j_3 = A_reg_bank58_p0_rd_data;	// matmul/matmul-hw.mlir:12273:32, :16188:5
  //PROBE: a_i_k_10_i_j_3	// matmul/matmul-hw.mlir:16189:5
  assign b_i_k_10_i_j_3 = _T_2617;	// matmul/matmul-hw.mlir:16191:5
  //PROBE: b_i_k_10_i_j_3	// matmul/matmul-hw.mlir:16192:5
  assign c_prev_i_k_10_i_j_3 = C_reg_bank10_p0_rd_data_2392;	// matmul/matmul-hw.mlir:15874:37, :16194:5
  //PROBE: c_prev_i_k_10_i_j_3	// matmul/matmul-hw.mlir:16195:5
  assign tk_i_k_10_i_j_3 = _T_2852;	// matmul/matmul-hw.mlir:16197:5
  //PROBE: tk_i_k_10_i_j_3	// matmul/matmul-hw.mlir:16198:5
  wire [31:0] _T_3172 = mult_inst58_result + C_reg_bank10_p0_rd_data_2392;	// matmul/matmul-hw.mlir:15874:37, :16185:27, :16199:13
  assign c_i_k_10_i_j_3 = _T_3172;	// matmul/matmul-hw.mlir:16201:5
  //PROBE: c_i_k_10_i_j_3	// matmul/matmul-hw.mlir:16202:5
  assign _T_1074 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16203:13
  assign _T_1073 = _T_2892 ? _T_3172 : 32'bx;	// matmul/matmul-hw.mlir:9108:19, :16204:13
  localparam [3:0] _T_3174 = 4'h0;	// matmul/matmul-hw.mlir:16207:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16208:5
    if (rst)	// matmul/matmul-hw.mlir:16208:5
      i_k_next_3173 <= _T_3174;	// matmul/matmul-hw.mlir:16211:7
    else	// matmul/matmul-hw.mlir:16208:5
      i_k_next_3173 <= i_k_next_3170;	// matmul/matmul-hw.mlir:16176:13, :16209:7
  end // always @(posedge)
  assign _T_1072 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16213:13
  assign _T_1071 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16214:13
  mult mult_inst59 (	// matmul/matmul-hw.mlir:16215:27
    .a      (A_reg_bank59_p0_rd_data),	// matmul/matmul-hw.mlir:12274:32
    .b      (_T_2633),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst59_result)
  );
  assign _T_1070 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16216:13
  assign a_i_k_11_i_j_3 = A_reg_bank59_p0_rd_data;	// matmul/matmul-hw.mlir:12274:32, :16218:5
  //PROBE: a_i_k_11_i_j_3	// matmul/matmul-hw.mlir:16219:5
  assign b_i_k_11_i_j_3 = _T_2633;	// matmul/matmul-hw.mlir:16221:5
  //PROBE: b_i_k_11_i_j_3	// matmul/matmul-hw.mlir:16222:5
  assign c_prev_i_k_11_i_j_3 = C_reg_bank11_p0_rd_data_2391;	// matmul/matmul-hw.mlir:15875:37, :16224:5
  //PROBE: c_prev_i_k_11_i_j_3	// matmul/matmul-hw.mlir:16225:5
  assign tk_i_k_11_i_j_3 = _T_2863;	// matmul/matmul-hw.mlir:16227:5
  //PROBE: tk_i_k_11_i_j_3	// matmul/matmul-hw.mlir:16228:5
  wire [31:0] _T_3175 = mult_inst59_result + C_reg_bank11_p0_rd_data_2391;	// matmul/matmul-hw.mlir:15875:37, :16215:27, :16229:13
  assign c_i_k_11_i_j_3 = _T_3175;	// matmul/matmul-hw.mlir:16231:5
  //PROBE: c_i_k_11_i_j_3	// matmul/matmul-hw.mlir:16232:5
  assign _T_1069 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16233:13
  assign _T_1068 = _T_2897 ? _T_3175 : 32'bx;	// matmul/matmul-hw.mlir:9103:19, :16234:13
  localparam [3:0] _T_3177 = 4'h0;	// matmul/matmul-hw.mlir:16237:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16238:5
    if (rst)	// matmul/matmul-hw.mlir:16238:5
      i_k_next_3176 <= _T_3177;	// matmul/matmul-hw.mlir:16241:7
    else	// matmul/matmul-hw.mlir:16238:5
      i_k_next_3176 <= i_k_next_3173;	// matmul/matmul-hw.mlir:16206:13, :16239:7
  end // always @(posedge)
  assign _T_1067 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16243:13
  assign _T_1066 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16244:13
  mult mult_inst60 (	// matmul/matmul-hw.mlir:16245:27
    .a      (A_reg_bank60_p0_rd_data),	// matmul/matmul-hw.mlir:12275:32
    .b      (_T_2649),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst60_result)
  );
  assign _T_1065 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16246:13
  assign a_i_k_12_i_j_3 = A_reg_bank60_p0_rd_data;	// matmul/matmul-hw.mlir:12275:32, :16248:5
  //PROBE: a_i_k_12_i_j_3	// matmul/matmul-hw.mlir:16249:5
  assign b_i_k_12_i_j_3 = _T_2649;	// matmul/matmul-hw.mlir:16251:5
  //PROBE: b_i_k_12_i_j_3	// matmul/matmul-hw.mlir:16252:5
  assign c_prev_i_k_12_i_j_3 = C_reg_bank12_p0_rd_data_2390;	// matmul/matmul-hw.mlir:15876:37, :16254:5
  //PROBE: c_prev_i_k_12_i_j_3	// matmul/matmul-hw.mlir:16255:5
  assign tk_i_k_12_i_j_3 = _T_2874;	// matmul/matmul-hw.mlir:16257:5
  //PROBE: tk_i_k_12_i_j_3	// matmul/matmul-hw.mlir:16258:5
  wire [31:0] _T_3178 = mult_inst60_result + C_reg_bank12_p0_rd_data_2390;	// matmul/matmul-hw.mlir:15876:37, :16245:27, :16259:13
  assign c_i_k_12_i_j_3 = _T_3178;	// matmul/matmul-hw.mlir:16261:5
  //PROBE: c_i_k_12_i_j_3	// matmul/matmul-hw.mlir:16262:5
  assign _T_1064 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16263:13
  assign _T_1063 = _T_2902 ? _T_3178 : 32'bx;	// matmul/matmul-hw.mlir:9098:19, :16264:13
  localparam [3:0] _T_3180 = 4'h0;	// matmul/matmul-hw.mlir:16267:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16268:5
    if (rst)	// matmul/matmul-hw.mlir:16268:5
      i_k_next_3179 <= _T_3180;	// matmul/matmul-hw.mlir:16271:7
    else	// matmul/matmul-hw.mlir:16268:5
      i_k_next_3179 <= i_k_next_3176;	// matmul/matmul-hw.mlir:16236:13, :16269:7
  end // always @(posedge)
  assign _T_1062 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16273:13
  assign _T_1061 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16274:13
  mult mult_inst61 (	// matmul/matmul-hw.mlir:16275:27
    .a      (A_reg_bank61_p0_rd_data),	// matmul/matmul-hw.mlir:12276:32
    .b      (_T_2665),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst61_result)
  );
  assign _T_1060 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16276:13
  assign a_i_k_13_i_j_3 = A_reg_bank61_p0_rd_data;	// matmul/matmul-hw.mlir:12276:32, :16278:5
  //PROBE: a_i_k_13_i_j_3	// matmul/matmul-hw.mlir:16279:5
  assign b_i_k_13_i_j_3 = _T_2665;	// matmul/matmul-hw.mlir:16281:5
  //PROBE: b_i_k_13_i_j_3	// matmul/matmul-hw.mlir:16282:5
  assign c_prev_i_k_13_i_j_3 = C_reg_bank13_p0_rd_data_2389;	// matmul/matmul-hw.mlir:15877:37, :16284:5
  //PROBE: c_prev_i_k_13_i_j_3	// matmul/matmul-hw.mlir:16285:5
  assign tk_i_k_13_i_j_3 = _T_2885;	// matmul/matmul-hw.mlir:16287:5
  //PROBE: tk_i_k_13_i_j_3	// matmul/matmul-hw.mlir:16288:5
  wire [31:0] _T_3181 = mult_inst61_result + C_reg_bank13_p0_rd_data_2389;	// matmul/matmul-hw.mlir:15877:37, :16275:27, :16289:13
  assign c_i_k_13_i_j_3 = _T_3181;	// matmul/matmul-hw.mlir:16291:5
  //PROBE: c_i_k_13_i_j_3	// matmul/matmul-hw.mlir:16292:5
  assign _T_1059 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16293:13
  assign _T_1058 = _T_2907 ? _T_3181 : 32'bx;	// matmul/matmul-hw.mlir:9093:19, :16294:13
  localparam [3:0] _T_3183 = 4'h0;	// matmul/matmul-hw.mlir:16297:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16298:5
    if (rst)	// matmul/matmul-hw.mlir:16298:5
      i_k_next_3182 <= _T_3183;	// matmul/matmul-hw.mlir:16301:7
    else	// matmul/matmul-hw.mlir:16298:5
      i_k_next_3182 <= i_k_next_3179;	// matmul/matmul-hw.mlir:16266:13, :16299:7
  end // always @(posedge)
  assign _T_1057 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16303:13
  assign _T_1056 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16304:13
  mult mult_inst62 (	// matmul/matmul-hw.mlir:16305:27
    .a      (A_reg_bank62_p0_rd_data),	// matmul/matmul-hw.mlir:12277:32
    .b      (_T_2681),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst62_result)
  );
  assign _T_1055 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16306:13
  assign a_i_k_14_i_j_3 = A_reg_bank62_p0_rd_data;	// matmul/matmul-hw.mlir:12277:32, :16308:5
  //PROBE: a_i_k_14_i_j_3	// matmul/matmul-hw.mlir:16309:5
  assign b_i_k_14_i_j_3 = _T_2681;	// matmul/matmul-hw.mlir:16311:5
  //PROBE: b_i_k_14_i_j_3	// matmul/matmul-hw.mlir:16312:5
  assign c_prev_i_k_14_i_j_3 = C_reg_bank14_p0_rd_data_2388;	// matmul/matmul-hw.mlir:15878:37, :16314:5
  //PROBE: c_prev_i_k_14_i_j_3	// matmul/matmul-hw.mlir:16315:5
  assign tk_i_k_14_i_j_3 = _T_2892;	// matmul/matmul-hw.mlir:16317:5
  //PROBE: tk_i_k_14_i_j_3	// matmul/matmul-hw.mlir:16318:5
  wire [31:0] _T_3184 = mult_inst62_result + C_reg_bank14_p0_rd_data_2388;	// matmul/matmul-hw.mlir:15878:37, :16305:27, :16319:13
  assign c_i_k_14_i_j_3 = _T_3184;	// matmul/matmul-hw.mlir:16321:5
  //PROBE: c_i_k_14_i_j_3	// matmul/matmul-hw.mlir:16322:5
  assign _T_1054 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16323:13
  assign _T_1053 = _T_2912 ? _T_3184 : 32'bx;	// matmul/matmul-hw.mlir:9088:19, :16324:13
  localparam [3:0] _T_3186 = 4'h0;	// matmul/matmul-hw.mlir:16327:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16328:5
    if (rst)	// matmul/matmul-hw.mlir:16328:5
      i_k_next_3185 <= _T_3186;	// matmul/matmul-hw.mlir:16331:7
    else	// matmul/matmul-hw.mlir:16328:5
      i_k_next_3185 <= i_k_next_3182;	// matmul/matmul-hw.mlir:16296:13, :16329:7
  end // always @(posedge)
  assign _T_1052 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16333:13
  assign _T_1051 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16334:13
  mult mult_inst63 (	// matmul/matmul-hw.mlir:16335:27
    .a      (A_reg_bank63_p0_rd_data),	// matmul/matmul-hw.mlir:12278:32
    .b      (_T_2697),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst63_result)
  );
  assign _T_1050 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16336:13
  assign a_i_k_15_i_j_3 = A_reg_bank63_p0_rd_data;	// matmul/matmul-hw.mlir:12278:32, :16338:5
  //PROBE: a_i_k_15_i_j_3	// matmul/matmul-hw.mlir:16339:5
  assign b_i_k_15_i_j_3 = _T_2697;	// matmul/matmul-hw.mlir:16341:5
  //PROBE: b_i_k_15_i_j_3	// matmul/matmul-hw.mlir:16342:5
  assign c_prev_i_k_15_i_j_3 = C_reg_bank15_p0_rd_data_2387;	// matmul/matmul-hw.mlir:15879:37, :16344:5
  //PROBE: c_prev_i_k_15_i_j_3	// matmul/matmul-hw.mlir:16345:5
  assign tk_i_k_15_i_j_3 = _T_2897;	// matmul/matmul-hw.mlir:16347:5
  //PROBE: tk_i_k_15_i_j_3	// matmul/matmul-hw.mlir:16348:5
  wire [31:0] _T_3187 = mult_inst63_result + C_reg_bank15_p0_rd_data_2387;	// matmul/matmul-hw.mlir:15879:37, :16335:27, :16349:13
  assign c_i_k_15_i_j_3 = _T_3187;	// matmul/matmul-hw.mlir:16351:5
  //PROBE: c_i_k_15_i_j_3	// matmul/matmul-hw.mlir:16352:5
  assign _T_1049 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16353:13
  assign _T_1048 = _T_2917 ? _T_3187 : 32'bx;	// matmul/matmul-hw.mlir:9083:19, :16354:13
  localparam [3:0] _T_3189 = 4'h0;	// matmul/matmul-hw.mlir:16357:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16358:5
    if (rst)	// matmul/matmul-hw.mlir:16358:5
      i_k_next_3188 <= _T_3189;	// matmul/matmul-hw.mlir:16361:7
    else	// matmul/matmul-hw.mlir:16358:5
      i_k_next_3188 <= i_k_next_3185;	// matmul/matmul-hw.mlir:16326:13, :16359:7
  end // always @(posedge)
  assign _T_1047 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16363:13
  wire [3:0][3:0] _T_3191 = i_delayed_3190;	// matmul/matmul-hw.mlir:16365:13
  wire [3:0][3:0] _T_3192 = {_T_3191[2'h0+:3], {{i_k_next_3188}}};	// matmul/matmul-hw.mlir:16356:13, :16366:19, :16367:13, :16368:13, :16369:13
  wire [3:0][3:0] _T_3193 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:16370:19, :16371:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16372:5
    if (rst)	// matmul/matmul-hw.mlir:16372:5
      i_delayed_3190 <= _T_3193;	// matmul/matmul-hw.mlir:16375:7
    else	// matmul/matmul-hw.mlir:16372:5
      i_delayed_3190 <= _T_3192;	// matmul/matmul-hw.mlir:16373:7
  end // always @(posedge)
  assign _T_1046 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16379:13
  assign _T_1045 = _T_2922 ? i_delayed_3190[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:9080:18, :16365:13, :16377:20, :16378:13, :16380:13
  assign _T_1044 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16381:13
  assign _T_1043 = _T_2922 ? C_reg_bank16_p0_rd_data_2386 : 32'bx;	// matmul/matmul-hw.mlir:9078:19, :15880:37, :16382:13
  localparam [3:0] _T_3195 = 4'h0;	// matmul/matmul-hw.mlir:16385:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16386:5
    if (rst)	// matmul/matmul-hw.mlir:16386:5
      i_j_next_3194 <= _T_3195;	// matmul/matmul-hw.mlir:16389:7
    else	// matmul/matmul-hw.mlir:16386:5
      i_j_next_3194 <= i_j_next_3123;	// matmul/matmul-hw.mlir:15789:13, :16387:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3196 (	// matmul/matmul-hw.mlir:16459:36
    .p0_rd_en   (_T_1038),	// matmul/matmul-hw.mlir:16481:13
    .p1_wr_en   (_T_1042),	// matmul/matmul-hw.mlir:16476:13
    .p1_wr_data (_T_1041),	// matmul/matmul-hw.mlir:16477:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2385)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3197 (	// matmul/matmul-hw.mlir:16460:36
    .p0_rd_en   (_T_1033),	// matmul/matmul-hw.mlir:16511:13
    .p1_wr_en   (_T_1037),	// matmul/matmul-hw.mlir:16498:13
    .p1_wr_data (_T_1036),	// matmul/matmul-hw.mlir:16499:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2384)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3198 (	// matmul/matmul-hw.mlir:16461:36
    .p0_rd_en   (_T_1028),	// matmul/matmul-hw.mlir:16541:13
    .p1_wr_en   (_T_1032),	// matmul/matmul-hw.mlir:16528:13
    .p1_wr_data (_T_1031),	// matmul/matmul-hw.mlir:16529:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2383)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3199 (	// matmul/matmul-hw.mlir:16462:36
    .p0_rd_en   (_T_1023),	// matmul/matmul-hw.mlir:16571:13
    .p1_wr_en   (_T_1027),	// matmul/matmul-hw.mlir:16558:13
    .p1_wr_data (_T_1026),	// matmul/matmul-hw.mlir:16559:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2382)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3200 (	// matmul/matmul-hw.mlir:16463:36
    .p0_rd_en   (_T_1018),	// matmul/matmul-hw.mlir:16601:13
    .p1_wr_en   (_T_1022),	// matmul/matmul-hw.mlir:16588:13
    .p1_wr_data (_T_1021),	// matmul/matmul-hw.mlir:16589:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2381)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3201 (	// matmul/matmul-hw.mlir:16464:36
    .p0_rd_en   (_T_1013),	// matmul/matmul-hw.mlir:16631:13
    .p1_wr_en   (_T_1017),	// matmul/matmul-hw.mlir:16618:13
    .p1_wr_data (_T_1016),	// matmul/matmul-hw.mlir:16619:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2380)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3202 (	// matmul/matmul-hw.mlir:16465:36
    .p0_rd_en   (_T_1008),	// matmul/matmul-hw.mlir:16661:13
    .p1_wr_en   (_T_1012),	// matmul/matmul-hw.mlir:16648:13
    .p1_wr_data (_T_1011),	// matmul/matmul-hw.mlir:16649:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2379)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3203 (	// matmul/matmul-hw.mlir:16466:36
    .p0_rd_en   (_T_1003),	// matmul/matmul-hw.mlir:16691:13
    .p1_wr_en   (_T_1007),	// matmul/matmul-hw.mlir:16678:13
    .p1_wr_data (_T_1006),	// matmul/matmul-hw.mlir:16679:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2378)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3204 (	// matmul/matmul-hw.mlir:16467:36
    .p0_rd_en   (_T_998),	// matmul/matmul-hw.mlir:16721:13
    .p1_wr_en   (_T_1002),	// matmul/matmul-hw.mlir:16708:13
    .p1_wr_data (_T_1001),	// matmul/matmul-hw.mlir:16709:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2377)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3205 (	// matmul/matmul-hw.mlir:16468:36
    .p0_rd_en   (_T_993),	// matmul/matmul-hw.mlir:16751:13
    .p1_wr_en   (_T_997),	// matmul/matmul-hw.mlir:16738:13
    .p1_wr_data (_T_996),	// matmul/matmul-hw.mlir:16739:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2376)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3206 (	// matmul/matmul-hw.mlir:16469:37
    .p0_rd_en   (_T_988),	// matmul/matmul-hw.mlir:16781:13
    .p1_wr_en   (_T_992),	// matmul/matmul-hw.mlir:16768:13
    .p1_wr_data (_T_991),	// matmul/matmul-hw.mlir:16769:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2375)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3207 (	// matmul/matmul-hw.mlir:16470:37
    .p0_rd_en   (_T_983),	// matmul/matmul-hw.mlir:16811:13
    .p1_wr_en   (_T_987),	// matmul/matmul-hw.mlir:16798:13
    .p1_wr_data (_T_986),	// matmul/matmul-hw.mlir:16799:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2374)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3208 (	// matmul/matmul-hw.mlir:16471:37
    .p0_rd_en   (_T_978),	// matmul/matmul-hw.mlir:16841:13
    .p1_wr_en   (_T_982),	// matmul/matmul-hw.mlir:16828:13
    .p1_wr_data (_T_981),	// matmul/matmul-hw.mlir:16829:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2373)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3209 (	// matmul/matmul-hw.mlir:16472:37
    .p0_rd_en   (_T_973),	// matmul/matmul-hw.mlir:16871:13
    .p1_wr_en   (_T_977),	// matmul/matmul-hw.mlir:16858:13
    .p1_wr_data (_T_976),	// matmul/matmul-hw.mlir:16859:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2372)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3210 (	// matmul/matmul-hw.mlir:16473:37
    .p0_rd_en   (_T_968),	// matmul/matmul-hw.mlir:16901:13
    .p1_wr_en   (_T_972),	// matmul/matmul-hw.mlir:16888:13
    .p1_wr_data (_T_971),	// matmul/matmul-hw.mlir:16889:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2371)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3211 (	// matmul/matmul-hw.mlir:16474:37
    .p0_rd_en   (_T_963),	// matmul/matmul-hw.mlir:16931:13
    .p1_wr_en   (_T_967),	// matmul/matmul-hw.mlir:16918:13
    .p1_wr_data (_T_966),	// matmul/matmul-hw.mlir:16919:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2370)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3212 (	// matmul/matmul-hw.mlir:16475:37
    .p0_rd_en   (_T_960),	// matmul/matmul-hw.mlir:16958:13
    .p1_wr_en   (_T_962),	// matmul/matmul-hw.mlir:16948:13
    .p1_wr_data (_T_961),	// matmul/matmul-hw.mlir:16949:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2369)
  );
  assign _T_1042 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16476:13
  assign _T_1041 = _T_2786 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :9076:19, :16477:13
  assign _T_1040 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16478:13
  assign _T_1039 = _T_2775 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16479:13
  mult mult_inst64 (	// matmul/matmul-hw.mlir:16480:27
    .a      (A_reg_bank64_p0_rd_data),	// matmul/matmul-hw.mlir:12279:32
    .b      (_T_2458),
    .t      (_T_2775),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst64_result)
  );
  assign _T_1038 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16481:13
  assign a_i_k_0_i_j_4 = A_reg_bank64_p0_rd_data;	// matmul/matmul-hw.mlir:12279:32, :16483:5
  //PROBE: a_i_k_0_i_j_4	// matmul/matmul-hw.mlir:16484:5
  assign b_i_k_0_i_j_4 = _T_2458;	// matmul/matmul-hw.mlir:16486:5
  //PROBE: b_i_k_0_i_j_4	// matmul/matmul-hw.mlir:16487:5
  assign c_prev_i_k_0_i_j_4 = C_reg_bank0_p0_rd_data_2385;	// matmul/matmul-hw.mlir:16459:36, :16489:5
  //PROBE: c_prev_i_k_0_i_j_4	// matmul/matmul-hw.mlir:16490:5
  assign tk_i_k_0_i_j_4 = _T_2753;	// matmul/matmul-hw.mlir:16492:5
  //PROBE: tk_i_k_0_i_j_4	// matmul/matmul-hw.mlir:16493:5
  wire [31:0] _T_3213 = mult_inst64_result + C_reg_bank0_p0_rd_data_2385;	// matmul/matmul-hw.mlir:16459:36, :16480:27, :16494:13
  assign c_i_k_0_i_j_4 = _T_3213;	// matmul/matmul-hw.mlir:16496:5
  //PROBE: c_i_k_0_i_j_4	// matmul/matmul-hw.mlir:16497:5
  assign _T_1037 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16498:13
  assign _T_1036 = _T_2797 ? _T_3213 : 32'bx;	// matmul/matmul-hw.mlir:9071:19, :16499:13
  localparam [3:0] _T_3215 = 4'h0;	// matmul/matmul-hw.mlir:16502:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16503:5
    if (rst)	// matmul/matmul-hw.mlir:16503:5
      i_k_next_3214 <= _T_3215;	// matmul/matmul-hw.mlir:16506:7
    else	// matmul/matmul-hw.mlir:16503:5
      i_k_next_3214 <= i_j_next_3194;	// matmul/matmul-hw.mlir:16384:13, :16504:7
  end // always @(posedge)
  assign _T_1035 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16508:13
  assign _T_1034 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16509:13
  mult mult_inst65 (	// matmul/matmul-hw.mlir:16510:27
    .a      (A_reg_bank65_p0_rd_data),	// matmul/matmul-hw.mlir:12280:32
    .b      (_T_2474),
    .t      (_T_2786),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst65_result)
  );
  assign _T_1033 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16511:13
  assign a_i_k_1_i_j_4 = A_reg_bank65_p0_rd_data;	// matmul/matmul-hw.mlir:12280:32, :16513:5
  //PROBE: a_i_k_1_i_j_4	// matmul/matmul-hw.mlir:16514:5
  assign b_i_k_1_i_j_4 = _T_2474;	// matmul/matmul-hw.mlir:16516:5
  //PROBE: b_i_k_1_i_j_4	// matmul/matmul-hw.mlir:16517:5
  assign c_prev_i_k_1_i_j_4 = C_reg_bank1_p0_rd_data_2384;	// matmul/matmul-hw.mlir:16460:36, :16519:5
  //PROBE: c_prev_i_k_1_i_j_4	// matmul/matmul-hw.mlir:16520:5
  assign tk_i_k_1_i_j_4 = _T_2764;	// matmul/matmul-hw.mlir:16522:5
  //PROBE: tk_i_k_1_i_j_4	// matmul/matmul-hw.mlir:16523:5
  wire [31:0] _T_3216 = mult_inst65_result + C_reg_bank1_p0_rd_data_2384;	// matmul/matmul-hw.mlir:16460:36, :16510:27, :16524:13
  assign c_i_k_1_i_j_4 = _T_3216;	// matmul/matmul-hw.mlir:16526:5
  //PROBE: c_i_k_1_i_j_4	// matmul/matmul-hw.mlir:16527:5
  assign _T_1032 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16528:13
  assign _T_1031 = _T_2808 ? _T_3216 : 32'bx;	// matmul/matmul-hw.mlir:9066:19, :16529:13
  localparam [3:0] _T_3218 = 4'h0;	// matmul/matmul-hw.mlir:16532:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16533:5
    if (rst)	// matmul/matmul-hw.mlir:16533:5
      i_k_next_3217 <= _T_3218;	// matmul/matmul-hw.mlir:16536:7
    else	// matmul/matmul-hw.mlir:16533:5
      i_k_next_3217 <= i_k_next_3214;	// matmul/matmul-hw.mlir:16501:13, :16534:7
  end // always @(posedge)
  assign _T_1030 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16538:13
  assign _T_1029 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16539:13
  mult mult_inst66 (	// matmul/matmul-hw.mlir:16540:27
    .a      (A_reg_bank66_p0_rd_data),	// matmul/matmul-hw.mlir:12281:32
    .b      (_T_2490),
    .t      (_T_2797),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst66_result)
  );
  assign _T_1028 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16541:13
  assign a_i_k_2_i_j_4 = A_reg_bank66_p0_rd_data;	// matmul/matmul-hw.mlir:12281:32, :16543:5
  //PROBE: a_i_k_2_i_j_4	// matmul/matmul-hw.mlir:16544:5
  assign b_i_k_2_i_j_4 = _T_2490;	// matmul/matmul-hw.mlir:16546:5
  //PROBE: b_i_k_2_i_j_4	// matmul/matmul-hw.mlir:16547:5
  assign c_prev_i_k_2_i_j_4 = C_reg_bank2_p0_rd_data_2383;	// matmul/matmul-hw.mlir:16461:36, :16549:5
  //PROBE: c_prev_i_k_2_i_j_4	// matmul/matmul-hw.mlir:16550:5
  assign tk_i_k_2_i_j_4 = _T_2775;	// matmul/matmul-hw.mlir:16552:5
  //PROBE: tk_i_k_2_i_j_4	// matmul/matmul-hw.mlir:16553:5
  wire [31:0] _T_3219 = mult_inst66_result + C_reg_bank2_p0_rd_data_2383;	// matmul/matmul-hw.mlir:16461:36, :16540:27, :16554:13
  assign c_i_k_2_i_j_4 = _T_3219;	// matmul/matmul-hw.mlir:16556:5
  //PROBE: c_i_k_2_i_j_4	// matmul/matmul-hw.mlir:16557:5
  assign _T_1027 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16558:13
  assign _T_1026 = _T_2819 ? _T_3219 : 32'bx;	// matmul/matmul-hw.mlir:9061:19, :16559:13
  localparam [3:0] _T_3221 = 4'h0;	// matmul/matmul-hw.mlir:16562:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16563:5
    if (rst)	// matmul/matmul-hw.mlir:16563:5
      i_k_next_3220 <= _T_3221;	// matmul/matmul-hw.mlir:16566:7
    else	// matmul/matmul-hw.mlir:16563:5
      i_k_next_3220 <= i_k_next_3217;	// matmul/matmul-hw.mlir:16531:13, :16564:7
  end // always @(posedge)
  assign _T_1025 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16568:13
  assign _T_1024 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16569:13
  mult mult_inst67 (	// matmul/matmul-hw.mlir:16570:27
    .a      (A_reg_bank67_p0_rd_data),	// matmul/matmul-hw.mlir:12282:32
    .b      (_T_2506),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst67_result)
  );
  assign _T_1023 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16571:13
  assign a_i_k_3_i_j_4 = A_reg_bank67_p0_rd_data;	// matmul/matmul-hw.mlir:12282:32, :16573:5
  //PROBE: a_i_k_3_i_j_4	// matmul/matmul-hw.mlir:16574:5
  assign b_i_k_3_i_j_4 = _T_2506;	// matmul/matmul-hw.mlir:16576:5
  //PROBE: b_i_k_3_i_j_4	// matmul/matmul-hw.mlir:16577:5
  assign c_prev_i_k_3_i_j_4 = C_reg_bank3_p0_rd_data_2382;	// matmul/matmul-hw.mlir:16462:36, :16579:5
  //PROBE: c_prev_i_k_3_i_j_4	// matmul/matmul-hw.mlir:16580:5
  assign tk_i_k_3_i_j_4 = _T_2786;	// matmul/matmul-hw.mlir:16582:5
  //PROBE: tk_i_k_3_i_j_4	// matmul/matmul-hw.mlir:16583:5
  wire [31:0] _T_3222 = mult_inst67_result + C_reg_bank3_p0_rd_data_2382;	// matmul/matmul-hw.mlir:16462:36, :16570:27, :16584:13
  assign c_i_k_3_i_j_4 = _T_3222;	// matmul/matmul-hw.mlir:16586:5
  //PROBE: c_i_k_3_i_j_4	// matmul/matmul-hw.mlir:16587:5
  assign _T_1022 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16588:13
  assign _T_1021 = _T_2830 ? _T_3222 : 32'bx;	// matmul/matmul-hw.mlir:9056:19, :16589:13
  localparam [3:0] _T_3224 = 4'h0;	// matmul/matmul-hw.mlir:16592:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16593:5
    if (rst)	// matmul/matmul-hw.mlir:16593:5
      i_k_next_3223 <= _T_3224;	// matmul/matmul-hw.mlir:16596:7
    else	// matmul/matmul-hw.mlir:16593:5
      i_k_next_3223 <= i_k_next_3220;	// matmul/matmul-hw.mlir:16561:13, :16594:7
  end // always @(posedge)
  assign _T_1020 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16598:13
  assign _T_1019 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16599:13
  mult mult_inst68 (	// matmul/matmul-hw.mlir:16600:27
    .a      (A_reg_bank68_p0_rd_data),	// matmul/matmul-hw.mlir:12283:32
    .b      (_T_2522),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst68_result)
  );
  assign _T_1018 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16601:13
  assign a_i_k_4_i_j_4 = A_reg_bank68_p0_rd_data;	// matmul/matmul-hw.mlir:12283:32, :16603:5
  //PROBE: a_i_k_4_i_j_4	// matmul/matmul-hw.mlir:16604:5
  assign b_i_k_4_i_j_4 = _T_2522;	// matmul/matmul-hw.mlir:16606:5
  //PROBE: b_i_k_4_i_j_4	// matmul/matmul-hw.mlir:16607:5
  assign c_prev_i_k_4_i_j_4 = C_reg_bank4_p0_rd_data_2381;	// matmul/matmul-hw.mlir:16463:36, :16609:5
  //PROBE: c_prev_i_k_4_i_j_4	// matmul/matmul-hw.mlir:16610:5
  assign tk_i_k_4_i_j_4 = _T_2797;	// matmul/matmul-hw.mlir:16612:5
  //PROBE: tk_i_k_4_i_j_4	// matmul/matmul-hw.mlir:16613:5
  wire [31:0] _T_3225 = mult_inst68_result + C_reg_bank4_p0_rd_data_2381;	// matmul/matmul-hw.mlir:16463:36, :16600:27, :16614:13
  assign c_i_k_4_i_j_4 = _T_3225;	// matmul/matmul-hw.mlir:16616:5
  //PROBE: c_i_k_4_i_j_4	// matmul/matmul-hw.mlir:16617:5
  assign _T_1017 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16618:13
  assign _T_1016 = _T_2841 ? _T_3225 : 32'bx;	// matmul/matmul-hw.mlir:9051:19, :16619:13
  localparam [3:0] _T_3227 = 4'h0;	// matmul/matmul-hw.mlir:16622:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16623:5
    if (rst)	// matmul/matmul-hw.mlir:16623:5
      i_k_next_3226 <= _T_3227;	// matmul/matmul-hw.mlir:16626:7
    else	// matmul/matmul-hw.mlir:16623:5
      i_k_next_3226 <= i_k_next_3223;	// matmul/matmul-hw.mlir:16591:13, :16624:7
  end // always @(posedge)
  assign _T_1015 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16628:13
  assign _T_1014 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16629:13
  mult mult_inst69 (	// matmul/matmul-hw.mlir:16630:27
    .a      (A_reg_bank69_p0_rd_data),	// matmul/matmul-hw.mlir:12284:32
    .b      (_T_2538),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst69_result)
  );
  assign _T_1013 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16631:13
  assign a_i_k_5_i_j_4 = A_reg_bank69_p0_rd_data;	// matmul/matmul-hw.mlir:12284:32, :16633:5
  //PROBE: a_i_k_5_i_j_4	// matmul/matmul-hw.mlir:16634:5
  assign b_i_k_5_i_j_4 = _T_2538;	// matmul/matmul-hw.mlir:16636:5
  //PROBE: b_i_k_5_i_j_4	// matmul/matmul-hw.mlir:16637:5
  assign c_prev_i_k_5_i_j_4 = C_reg_bank5_p0_rd_data_2380;	// matmul/matmul-hw.mlir:16464:36, :16639:5
  //PROBE: c_prev_i_k_5_i_j_4	// matmul/matmul-hw.mlir:16640:5
  assign tk_i_k_5_i_j_4 = _T_2808;	// matmul/matmul-hw.mlir:16642:5
  //PROBE: tk_i_k_5_i_j_4	// matmul/matmul-hw.mlir:16643:5
  wire [31:0] _T_3228 = mult_inst69_result + C_reg_bank5_p0_rd_data_2380;	// matmul/matmul-hw.mlir:16464:36, :16630:27, :16644:13
  assign c_i_k_5_i_j_4 = _T_3228;	// matmul/matmul-hw.mlir:16646:5
  //PROBE: c_i_k_5_i_j_4	// matmul/matmul-hw.mlir:16647:5
  assign _T_1012 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16648:13
  assign _T_1011 = _T_2852 ? _T_3228 : 32'bx;	// matmul/matmul-hw.mlir:9046:19, :16649:13
  localparam [3:0] _T_3230 = 4'h0;	// matmul/matmul-hw.mlir:16652:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16653:5
    if (rst)	// matmul/matmul-hw.mlir:16653:5
      i_k_next_3229 <= _T_3230;	// matmul/matmul-hw.mlir:16656:7
    else	// matmul/matmul-hw.mlir:16653:5
      i_k_next_3229 <= i_k_next_3226;	// matmul/matmul-hw.mlir:16621:13, :16654:7
  end // always @(posedge)
  assign _T_1010 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16658:13
  assign _T_1009 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16659:13
  mult mult_inst70 (	// matmul/matmul-hw.mlir:16660:27
    .a      (A_reg_bank70_p0_rd_data),	// matmul/matmul-hw.mlir:12285:32
    .b      (_T_2554),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst70_result)
  );
  assign _T_1008 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16661:13
  assign a_i_k_6_i_j_4 = A_reg_bank70_p0_rd_data;	// matmul/matmul-hw.mlir:12285:32, :16663:5
  //PROBE: a_i_k_6_i_j_4	// matmul/matmul-hw.mlir:16664:5
  assign b_i_k_6_i_j_4 = _T_2554;	// matmul/matmul-hw.mlir:16666:5
  //PROBE: b_i_k_6_i_j_4	// matmul/matmul-hw.mlir:16667:5
  assign c_prev_i_k_6_i_j_4 = C_reg_bank6_p0_rd_data_2379;	// matmul/matmul-hw.mlir:16465:36, :16669:5
  //PROBE: c_prev_i_k_6_i_j_4	// matmul/matmul-hw.mlir:16670:5
  assign tk_i_k_6_i_j_4 = _T_2819;	// matmul/matmul-hw.mlir:16672:5
  //PROBE: tk_i_k_6_i_j_4	// matmul/matmul-hw.mlir:16673:5
  wire [31:0] _T_3231 = mult_inst70_result + C_reg_bank6_p0_rd_data_2379;	// matmul/matmul-hw.mlir:16465:36, :16660:27, :16674:13
  assign c_i_k_6_i_j_4 = _T_3231;	// matmul/matmul-hw.mlir:16676:5
  //PROBE: c_i_k_6_i_j_4	// matmul/matmul-hw.mlir:16677:5
  assign _T_1007 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16678:13
  assign _T_1006 = _T_2863 ? _T_3231 : 32'bx;	// matmul/matmul-hw.mlir:9041:19, :16679:13
  localparam [3:0] _T_3233 = 4'h0;	// matmul/matmul-hw.mlir:16682:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16683:5
    if (rst)	// matmul/matmul-hw.mlir:16683:5
      i_k_next_3232 <= _T_3233;	// matmul/matmul-hw.mlir:16686:7
    else	// matmul/matmul-hw.mlir:16683:5
      i_k_next_3232 <= i_k_next_3229;	// matmul/matmul-hw.mlir:16651:13, :16684:7
  end // always @(posedge)
  assign _T_1005 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16688:13
  assign _T_1004 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16689:13
  mult mult_inst71 (	// matmul/matmul-hw.mlir:16690:27
    .a      (A_reg_bank71_p0_rd_data),	// matmul/matmul-hw.mlir:12286:32
    .b      (_T_2570),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst71_result)
  );
  assign _T_1003 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16691:13
  assign a_i_k_7_i_j_4 = A_reg_bank71_p0_rd_data;	// matmul/matmul-hw.mlir:12286:32, :16693:5
  //PROBE: a_i_k_7_i_j_4	// matmul/matmul-hw.mlir:16694:5
  assign b_i_k_7_i_j_4 = _T_2570;	// matmul/matmul-hw.mlir:16696:5
  //PROBE: b_i_k_7_i_j_4	// matmul/matmul-hw.mlir:16697:5
  assign c_prev_i_k_7_i_j_4 = C_reg_bank7_p0_rd_data_2378;	// matmul/matmul-hw.mlir:16466:36, :16699:5
  //PROBE: c_prev_i_k_7_i_j_4	// matmul/matmul-hw.mlir:16700:5
  assign tk_i_k_7_i_j_4 = _T_2830;	// matmul/matmul-hw.mlir:16702:5
  //PROBE: tk_i_k_7_i_j_4	// matmul/matmul-hw.mlir:16703:5
  wire [31:0] _T_3234 = mult_inst71_result + C_reg_bank7_p0_rd_data_2378;	// matmul/matmul-hw.mlir:16466:36, :16690:27, :16704:13
  assign c_i_k_7_i_j_4 = _T_3234;	// matmul/matmul-hw.mlir:16706:5
  //PROBE: c_i_k_7_i_j_4	// matmul/matmul-hw.mlir:16707:5
  assign _T_1002 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16708:13
  assign _T_1001 = _T_2874 ? _T_3234 : 32'bx;	// matmul/matmul-hw.mlir:9036:19, :16709:13
  localparam [3:0] _T_3236 = 4'h0;	// matmul/matmul-hw.mlir:16712:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16713:5
    if (rst)	// matmul/matmul-hw.mlir:16713:5
      i_k_next_3235 <= _T_3236;	// matmul/matmul-hw.mlir:16716:7
    else	// matmul/matmul-hw.mlir:16713:5
      i_k_next_3235 <= i_k_next_3232;	// matmul/matmul-hw.mlir:16681:13, :16714:7
  end // always @(posedge)
  assign _T_1000 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16718:13
  assign _T_999 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16719:13
  mult mult_inst72 (	// matmul/matmul-hw.mlir:16720:27
    .a      (A_reg_bank72_p0_rd_data),	// matmul/matmul-hw.mlir:12287:32
    .b      (_T_2586),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst72_result)
  );
  assign _T_998 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16721:13
  assign a_i_k_8_i_j_4 = A_reg_bank72_p0_rd_data;	// matmul/matmul-hw.mlir:12287:32, :16723:5
  //PROBE: a_i_k_8_i_j_4	// matmul/matmul-hw.mlir:16724:5
  assign b_i_k_8_i_j_4 = _T_2586;	// matmul/matmul-hw.mlir:16726:5
  //PROBE: b_i_k_8_i_j_4	// matmul/matmul-hw.mlir:16727:5
  assign c_prev_i_k_8_i_j_4 = C_reg_bank8_p0_rd_data_2377;	// matmul/matmul-hw.mlir:16467:36, :16729:5
  //PROBE: c_prev_i_k_8_i_j_4	// matmul/matmul-hw.mlir:16730:5
  assign tk_i_k_8_i_j_4 = _T_2841;	// matmul/matmul-hw.mlir:16732:5
  //PROBE: tk_i_k_8_i_j_4	// matmul/matmul-hw.mlir:16733:5
  wire [31:0] _T_3237 = mult_inst72_result + C_reg_bank8_p0_rd_data_2377;	// matmul/matmul-hw.mlir:16467:36, :16720:27, :16734:13
  assign c_i_k_8_i_j_4 = _T_3237;	// matmul/matmul-hw.mlir:16736:5
  //PROBE: c_i_k_8_i_j_4	// matmul/matmul-hw.mlir:16737:5
  assign _T_997 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16738:13
  assign _T_996 = _T_2885 ? _T_3237 : 32'bx;	// matmul/matmul-hw.mlir:9031:19, :16739:13
  localparam [3:0] _T_3239 = 4'h0;	// matmul/matmul-hw.mlir:16742:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16743:5
    if (rst)	// matmul/matmul-hw.mlir:16743:5
      i_k_next_3238 <= _T_3239;	// matmul/matmul-hw.mlir:16746:7
    else	// matmul/matmul-hw.mlir:16743:5
      i_k_next_3238 <= i_k_next_3235;	// matmul/matmul-hw.mlir:16711:13, :16744:7
  end // always @(posedge)
  assign _T_995 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16748:13
  assign _T_994 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16749:13
  mult mult_inst73 (	// matmul/matmul-hw.mlir:16750:27
    .a      (A_reg_bank73_p0_rd_data),	// matmul/matmul-hw.mlir:12288:32
    .b      (_T_2602),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst73_result)
  );
  assign _T_993 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16751:13
  assign a_i_k_9_i_j_4 = A_reg_bank73_p0_rd_data;	// matmul/matmul-hw.mlir:12288:32, :16753:5
  //PROBE: a_i_k_9_i_j_4	// matmul/matmul-hw.mlir:16754:5
  assign b_i_k_9_i_j_4 = _T_2602;	// matmul/matmul-hw.mlir:16756:5
  //PROBE: b_i_k_9_i_j_4	// matmul/matmul-hw.mlir:16757:5
  assign c_prev_i_k_9_i_j_4 = C_reg_bank9_p0_rd_data_2376;	// matmul/matmul-hw.mlir:16468:36, :16759:5
  //PROBE: c_prev_i_k_9_i_j_4	// matmul/matmul-hw.mlir:16760:5
  assign tk_i_k_9_i_j_4 = _T_2852;	// matmul/matmul-hw.mlir:16762:5
  //PROBE: tk_i_k_9_i_j_4	// matmul/matmul-hw.mlir:16763:5
  wire [31:0] _T_3240 = mult_inst73_result + C_reg_bank9_p0_rd_data_2376;	// matmul/matmul-hw.mlir:16468:36, :16750:27, :16764:13
  assign c_i_k_9_i_j_4 = _T_3240;	// matmul/matmul-hw.mlir:16766:5
  //PROBE: c_i_k_9_i_j_4	// matmul/matmul-hw.mlir:16767:5
  assign _T_992 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16768:13
  assign _T_991 = _T_2892 ? _T_3240 : 32'bx;	// matmul/matmul-hw.mlir:9026:19, :16769:13
  localparam [3:0] _T_3242 = 4'h0;	// matmul/matmul-hw.mlir:16772:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16773:5
    if (rst)	// matmul/matmul-hw.mlir:16773:5
      i_k_next_3241 <= _T_3242;	// matmul/matmul-hw.mlir:16776:7
    else	// matmul/matmul-hw.mlir:16773:5
      i_k_next_3241 <= i_k_next_3238;	// matmul/matmul-hw.mlir:16741:13, :16774:7
  end // always @(posedge)
  assign _T_990 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16778:13
  assign _T_989 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16779:13
  mult mult_inst74 (	// matmul/matmul-hw.mlir:16780:27
    .a      (A_reg_bank74_p0_rd_data),	// matmul/matmul-hw.mlir:12289:32
    .b      (_T_2618),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst74_result)
  );
  assign _T_988 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16781:13
  assign a_i_k_10_i_j_4 = A_reg_bank74_p0_rd_data;	// matmul/matmul-hw.mlir:12289:32, :16783:5
  //PROBE: a_i_k_10_i_j_4	// matmul/matmul-hw.mlir:16784:5
  assign b_i_k_10_i_j_4 = _T_2618;	// matmul/matmul-hw.mlir:16786:5
  //PROBE: b_i_k_10_i_j_4	// matmul/matmul-hw.mlir:16787:5
  assign c_prev_i_k_10_i_j_4 = C_reg_bank10_p0_rd_data_2375;	// matmul/matmul-hw.mlir:16469:37, :16789:5
  //PROBE: c_prev_i_k_10_i_j_4	// matmul/matmul-hw.mlir:16790:5
  assign tk_i_k_10_i_j_4 = _T_2863;	// matmul/matmul-hw.mlir:16792:5
  //PROBE: tk_i_k_10_i_j_4	// matmul/matmul-hw.mlir:16793:5
  wire [31:0] _T_3243 = mult_inst74_result + C_reg_bank10_p0_rd_data_2375;	// matmul/matmul-hw.mlir:16469:37, :16780:27, :16794:13
  assign c_i_k_10_i_j_4 = _T_3243;	// matmul/matmul-hw.mlir:16796:5
  //PROBE: c_i_k_10_i_j_4	// matmul/matmul-hw.mlir:16797:5
  assign _T_987 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16798:13
  assign _T_986 = _T_2897 ? _T_3243 : 32'bx;	// matmul/matmul-hw.mlir:9021:19, :16799:13
  localparam [3:0] _T_3245 = 4'h0;	// matmul/matmul-hw.mlir:16802:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16803:5
    if (rst)	// matmul/matmul-hw.mlir:16803:5
      i_k_next_3244 <= _T_3245;	// matmul/matmul-hw.mlir:16806:7
    else	// matmul/matmul-hw.mlir:16803:5
      i_k_next_3244 <= i_k_next_3241;	// matmul/matmul-hw.mlir:16771:13, :16804:7
  end // always @(posedge)
  assign _T_985 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16808:13
  assign _T_984 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16809:13
  mult mult_inst75 (	// matmul/matmul-hw.mlir:16810:27
    .a      (A_reg_bank75_p0_rd_data),	// matmul/matmul-hw.mlir:12290:32
    .b      (_T_2634),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst75_result)
  );
  assign _T_983 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16811:13
  assign a_i_k_11_i_j_4 = A_reg_bank75_p0_rd_data;	// matmul/matmul-hw.mlir:12290:32, :16813:5
  //PROBE: a_i_k_11_i_j_4	// matmul/matmul-hw.mlir:16814:5
  assign b_i_k_11_i_j_4 = _T_2634;	// matmul/matmul-hw.mlir:16816:5
  //PROBE: b_i_k_11_i_j_4	// matmul/matmul-hw.mlir:16817:5
  assign c_prev_i_k_11_i_j_4 = C_reg_bank11_p0_rd_data_2374;	// matmul/matmul-hw.mlir:16470:37, :16819:5
  //PROBE: c_prev_i_k_11_i_j_4	// matmul/matmul-hw.mlir:16820:5
  assign tk_i_k_11_i_j_4 = _T_2874;	// matmul/matmul-hw.mlir:16822:5
  //PROBE: tk_i_k_11_i_j_4	// matmul/matmul-hw.mlir:16823:5
  wire [31:0] _T_3246 = mult_inst75_result + C_reg_bank11_p0_rd_data_2374;	// matmul/matmul-hw.mlir:16470:37, :16810:27, :16824:13
  assign c_i_k_11_i_j_4 = _T_3246;	// matmul/matmul-hw.mlir:16826:5
  //PROBE: c_i_k_11_i_j_4	// matmul/matmul-hw.mlir:16827:5
  assign _T_982 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16828:13
  assign _T_981 = _T_2902 ? _T_3246 : 32'bx;	// matmul/matmul-hw.mlir:9016:19, :16829:13
  localparam [3:0] _T_3248 = 4'h0;	// matmul/matmul-hw.mlir:16832:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16833:5
    if (rst)	// matmul/matmul-hw.mlir:16833:5
      i_k_next_3247 <= _T_3248;	// matmul/matmul-hw.mlir:16836:7
    else	// matmul/matmul-hw.mlir:16833:5
      i_k_next_3247 <= i_k_next_3244;	// matmul/matmul-hw.mlir:16801:13, :16834:7
  end // always @(posedge)
  assign _T_980 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16838:13
  assign _T_979 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16839:13
  mult mult_inst76 (	// matmul/matmul-hw.mlir:16840:27
    .a      (A_reg_bank76_p0_rd_data),	// matmul/matmul-hw.mlir:12291:32
    .b      (_T_2650),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst76_result)
  );
  assign _T_978 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16841:13
  assign a_i_k_12_i_j_4 = A_reg_bank76_p0_rd_data;	// matmul/matmul-hw.mlir:12291:32, :16843:5
  //PROBE: a_i_k_12_i_j_4	// matmul/matmul-hw.mlir:16844:5
  assign b_i_k_12_i_j_4 = _T_2650;	// matmul/matmul-hw.mlir:16846:5
  //PROBE: b_i_k_12_i_j_4	// matmul/matmul-hw.mlir:16847:5
  assign c_prev_i_k_12_i_j_4 = C_reg_bank12_p0_rd_data_2373;	// matmul/matmul-hw.mlir:16471:37, :16849:5
  //PROBE: c_prev_i_k_12_i_j_4	// matmul/matmul-hw.mlir:16850:5
  assign tk_i_k_12_i_j_4 = _T_2885;	// matmul/matmul-hw.mlir:16852:5
  //PROBE: tk_i_k_12_i_j_4	// matmul/matmul-hw.mlir:16853:5
  wire [31:0] _T_3249 = mult_inst76_result + C_reg_bank12_p0_rd_data_2373;	// matmul/matmul-hw.mlir:16471:37, :16840:27, :16854:13
  assign c_i_k_12_i_j_4 = _T_3249;	// matmul/matmul-hw.mlir:16856:5
  //PROBE: c_i_k_12_i_j_4	// matmul/matmul-hw.mlir:16857:5
  assign _T_977 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16858:13
  assign _T_976 = _T_2907 ? _T_3249 : 32'bx;	// matmul/matmul-hw.mlir:9011:19, :16859:13
  localparam [3:0] _T_3251 = 4'h0;	// matmul/matmul-hw.mlir:16862:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16863:5
    if (rst)	// matmul/matmul-hw.mlir:16863:5
      i_k_next_3250 <= _T_3251;	// matmul/matmul-hw.mlir:16866:7
    else	// matmul/matmul-hw.mlir:16863:5
      i_k_next_3250 <= i_k_next_3247;	// matmul/matmul-hw.mlir:16831:13, :16864:7
  end // always @(posedge)
  assign _T_975 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16868:13
  assign _T_974 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16869:13
  mult mult_inst77 (	// matmul/matmul-hw.mlir:16870:27
    .a      (A_reg_bank77_p0_rd_data),	// matmul/matmul-hw.mlir:12292:32
    .b      (_T_2666),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst77_result)
  );
  assign _T_973 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16871:13
  assign a_i_k_13_i_j_4 = A_reg_bank77_p0_rd_data;	// matmul/matmul-hw.mlir:12292:32, :16873:5
  //PROBE: a_i_k_13_i_j_4	// matmul/matmul-hw.mlir:16874:5
  assign b_i_k_13_i_j_4 = _T_2666;	// matmul/matmul-hw.mlir:16876:5
  //PROBE: b_i_k_13_i_j_4	// matmul/matmul-hw.mlir:16877:5
  assign c_prev_i_k_13_i_j_4 = C_reg_bank13_p0_rd_data_2372;	// matmul/matmul-hw.mlir:16472:37, :16879:5
  //PROBE: c_prev_i_k_13_i_j_4	// matmul/matmul-hw.mlir:16880:5
  assign tk_i_k_13_i_j_4 = _T_2892;	// matmul/matmul-hw.mlir:16882:5
  //PROBE: tk_i_k_13_i_j_4	// matmul/matmul-hw.mlir:16883:5
  wire [31:0] _T_3252 = mult_inst77_result + C_reg_bank13_p0_rd_data_2372;	// matmul/matmul-hw.mlir:16472:37, :16870:27, :16884:13
  assign c_i_k_13_i_j_4 = _T_3252;	// matmul/matmul-hw.mlir:16886:5
  //PROBE: c_i_k_13_i_j_4	// matmul/matmul-hw.mlir:16887:5
  assign _T_972 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16888:13
  assign _T_971 = _T_2912 ? _T_3252 : 32'bx;	// matmul/matmul-hw.mlir:9006:19, :16889:13
  localparam [3:0] _T_3254 = 4'h0;	// matmul/matmul-hw.mlir:16892:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16893:5
    if (rst)	// matmul/matmul-hw.mlir:16893:5
      i_k_next_3253 <= _T_3254;	// matmul/matmul-hw.mlir:16896:7
    else	// matmul/matmul-hw.mlir:16893:5
      i_k_next_3253 <= i_k_next_3250;	// matmul/matmul-hw.mlir:16861:13, :16894:7
  end // always @(posedge)
  assign _T_970 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16898:13
  assign _T_969 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16899:13
  mult mult_inst78 (	// matmul/matmul-hw.mlir:16900:27
    .a      (A_reg_bank78_p0_rd_data),	// matmul/matmul-hw.mlir:12293:32
    .b      (_T_2682),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst78_result)
  );
  assign _T_968 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16901:13
  assign a_i_k_14_i_j_4 = A_reg_bank78_p0_rd_data;	// matmul/matmul-hw.mlir:12293:32, :16903:5
  //PROBE: a_i_k_14_i_j_4	// matmul/matmul-hw.mlir:16904:5
  assign b_i_k_14_i_j_4 = _T_2682;	// matmul/matmul-hw.mlir:16906:5
  //PROBE: b_i_k_14_i_j_4	// matmul/matmul-hw.mlir:16907:5
  assign c_prev_i_k_14_i_j_4 = C_reg_bank14_p0_rd_data_2371;	// matmul/matmul-hw.mlir:16473:37, :16909:5
  //PROBE: c_prev_i_k_14_i_j_4	// matmul/matmul-hw.mlir:16910:5
  assign tk_i_k_14_i_j_4 = _T_2897;	// matmul/matmul-hw.mlir:16912:5
  //PROBE: tk_i_k_14_i_j_4	// matmul/matmul-hw.mlir:16913:5
  wire [31:0] _T_3255 = mult_inst78_result + C_reg_bank14_p0_rd_data_2371;	// matmul/matmul-hw.mlir:16473:37, :16900:27, :16914:13
  assign c_i_k_14_i_j_4 = _T_3255;	// matmul/matmul-hw.mlir:16916:5
  //PROBE: c_i_k_14_i_j_4	// matmul/matmul-hw.mlir:16917:5
  assign _T_967 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16918:13
  assign _T_966 = _T_2917 ? _T_3255 : 32'bx;	// matmul/matmul-hw.mlir:9001:19, :16919:13
  localparam [3:0] _T_3257 = 4'h0;	// matmul/matmul-hw.mlir:16922:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16923:5
    if (rst)	// matmul/matmul-hw.mlir:16923:5
      i_k_next_3256 <= _T_3257;	// matmul/matmul-hw.mlir:16926:7
    else	// matmul/matmul-hw.mlir:16923:5
      i_k_next_3256 <= i_k_next_3253;	// matmul/matmul-hw.mlir:16891:13, :16924:7
  end // always @(posedge)
  assign _T_965 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16928:13
  assign _T_964 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16929:13
  mult mult_inst79 (	// matmul/matmul-hw.mlir:16930:27
    .a      (A_reg_bank79_p0_rd_data),	// matmul/matmul-hw.mlir:12294:32
    .b      (_T_2698),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst79_result)
  );
  assign _T_963 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16931:13
  assign a_i_k_15_i_j_4 = A_reg_bank79_p0_rd_data;	// matmul/matmul-hw.mlir:12294:32, :16933:5
  //PROBE: a_i_k_15_i_j_4	// matmul/matmul-hw.mlir:16934:5
  assign b_i_k_15_i_j_4 = _T_2698;	// matmul/matmul-hw.mlir:16936:5
  //PROBE: b_i_k_15_i_j_4	// matmul/matmul-hw.mlir:16937:5
  assign c_prev_i_k_15_i_j_4 = C_reg_bank15_p0_rd_data_2370;	// matmul/matmul-hw.mlir:16474:37, :16939:5
  //PROBE: c_prev_i_k_15_i_j_4	// matmul/matmul-hw.mlir:16940:5
  assign tk_i_k_15_i_j_4 = _T_2902;	// matmul/matmul-hw.mlir:16942:5
  //PROBE: tk_i_k_15_i_j_4	// matmul/matmul-hw.mlir:16943:5
  wire [31:0] _T_3258 = mult_inst79_result + C_reg_bank15_p0_rd_data_2370;	// matmul/matmul-hw.mlir:16474:37, :16930:27, :16944:13
  assign c_i_k_15_i_j_4 = _T_3258;	// matmul/matmul-hw.mlir:16946:5
  //PROBE: c_i_k_15_i_j_4	// matmul/matmul-hw.mlir:16947:5
  assign _T_962 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16948:13
  assign _T_961 = _T_2922 ? _T_3258 : 32'bx;	// matmul/matmul-hw.mlir:8996:19, :16949:13
  localparam [3:0] _T_3260 = 4'h0;	// matmul/matmul-hw.mlir:16952:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16953:5
    if (rst)	// matmul/matmul-hw.mlir:16953:5
      i_k_next_3259 <= _T_3260;	// matmul/matmul-hw.mlir:16956:7
    else	// matmul/matmul-hw.mlir:16953:5
      i_k_next_3259 <= i_k_next_3256;	// matmul/matmul-hw.mlir:16921:13, :16954:7
  end // always @(posedge)
  assign _T_960 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16958:13
  wire [3:0][3:0] _T_3262 = i_delayed_3261;	// matmul/matmul-hw.mlir:16960:13
  wire [3:0][3:0] _T_3263 = {_T_3262[2'h0+:3], {{i_k_next_3259}}};	// matmul/matmul-hw.mlir:16951:13, :16961:19, :16962:13, :16963:13, :16964:13
  wire [3:0][3:0] _T_3264 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:16965:19, :16966:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16967:5
    if (rst)	// matmul/matmul-hw.mlir:16967:5
      i_delayed_3261 <= _T_3264;	// matmul/matmul-hw.mlir:16970:7
    else	// matmul/matmul-hw.mlir:16967:5
      i_delayed_3261 <= _T_3263;	// matmul/matmul-hw.mlir:16968:7
  end // always @(posedge)
  assign _T_959 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16974:13
  assign _T_958 = _T_2927 ? i_delayed_3261[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8993:18, :16960:13, :16972:20, :16973:13, :16975:13
  assign _T_957 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :16976:13
  assign _T_956 = _T_2927 ? C_reg_bank16_p0_rd_data_2369 : 32'bx;	// matmul/matmul-hw.mlir:8991:19, :16475:37, :16977:13
  localparam [3:0] _T_3266 = 4'h0;	// matmul/matmul-hw.mlir:16980:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:16981:5
    if (rst)	// matmul/matmul-hw.mlir:16981:5
      i_j_next_3265 <= _T_3266;	// matmul/matmul-hw.mlir:16984:7
    else	// matmul/matmul-hw.mlir:16981:5
      i_j_next_3265 <= i_j_next_3194;	// matmul/matmul-hw.mlir:16384:13, :16982:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3267 (	// matmul/matmul-hw.mlir:17054:36
    .p0_rd_en   (_T_951),	// matmul/matmul-hw.mlir:17076:13
    .p1_wr_en   (_T_955),	// matmul/matmul-hw.mlir:17071:13
    .p1_wr_data (_T_954),	// matmul/matmul-hw.mlir:17072:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2368)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3268 (	// matmul/matmul-hw.mlir:17055:36
    .p0_rd_en   (_T_946),	// matmul/matmul-hw.mlir:17106:13
    .p1_wr_en   (_T_950),	// matmul/matmul-hw.mlir:17093:13
    .p1_wr_data (_T_949),	// matmul/matmul-hw.mlir:17094:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2367)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3269 (	// matmul/matmul-hw.mlir:17056:36
    .p0_rd_en   (_T_941),	// matmul/matmul-hw.mlir:17136:13
    .p1_wr_en   (_T_945),	// matmul/matmul-hw.mlir:17123:13
    .p1_wr_data (_T_944),	// matmul/matmul-hw.mlir:17124:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2366)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3270 (	// matmul/matmul-hw.mlir:17057:36
    .p0_rd_en   (_T_936),	// matmul/matmul-hw.mlir:17166:13
    .p1_wr_en   (_T_940),	// matmul/matmul-hw.mlir:17153:13
    .p1_wr_data (_T_939),	// matmul/matmul-hw.mlir:17154:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2365)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3271 (	// matmul/matmul-hw.mlir:17058:36
    .p0_rd_en   (_T_931),	// matmul/matmul-hw.mlir:17196:13
    .p1_wr_en   (_T_935),	// matmul/matmul-hw.mlir:17183:13
    .p1_wr_data (_T_934),	// matmul/matmul-hw.mlir:17184:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2364)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3272 (	// matmul/matmul-hw.mlir:17059:36
    .p0_rd_en   (_T_926),	// matmul/matmul-hw.mlir:17226:13
    .p1_wr_en   (_T_930),	// matmul/matmul-hw.mlir:17213:13
    .p1_wr_data (_T_929),	// matmul/matmul-hw.mlir:17214:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2363)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3273 (	// matmul/matmul-hw.mlir:17060:36
    .p0_rd_en   (_T_921),	// matmul/matmul-hw.mlir:17256:13
    .p1_wr_en   (_T_925),	// matmul/matmul-hw.mlir:17243:13
    .p1_wr_data (_T_924),	// matmul/matmul-hw.mlir:17244:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2362)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3274 (	// matmul/matmul-hw.mlir:17061:36
    .p0_rd_en   (_T_916),	// matmul/matmul-hw.mlir:17286:13
    .p1_wr_en   (_T_920),	// matmul/matmul-hw.mlir:17273:13
    .p1_wr_data (_T_919),	// matmul/matmul-hw.mlir:17274:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2361)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3275 (	// matmul/matmul-hw.mlir:17062:36
    .p0_rd_en   (_T_911),	// matmul/matmul-hw.mlir:17316:13
    .p1_wr_en   (_T_915),	// matmul/matmul-hw.mlir:17303:13
    .p1_wr_data (_T_914),	// matmul/matmul-hw.mlir:17304:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2360)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3276 (	// matmul/matmul-hw.mlir:17063:36
    .p0_rd_en   (_T_906),	// matmul/matmul-hw.mlir:17346:13
    .p1_wr_en   (_T_910),	// matmul/matmul-hw.mlir:17333:13
    .p1_wr_data (_T_909),	// matmul/matmul-hw.mlir:17334:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2359)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3277 (	// matmul/matmul-hw.mlir:17064:37
    .p0_rd_en   (_T_901),	// matmul/matmul-hw.mlir:17376:13
    .p1_wr_en   (_T_905),	// matmul/matmul-hw.mlir:17363:13
    .p1_wr_data (_T_904),	// matmul/matmul-hw.mlir:17364:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2358)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3278 (	// matmul/matmul-hw.mlir:17065:37
    .p0_rd_en   (_T_896),	// matmul/matmul-hw.mlir:17406:13
    .p1_wr_en   (_T_900),	// matmul/matmul-hw.mlir:17393:13
    .p1_wr_data (_T_899),	// matmul/matmul-hw.mlir:17394:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2357)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3279 (	// matmul/matmul-hw.mlir:17066:37
    .p0_rd_en   (_T_891),	// matmul/matmul-hw.mlir:17436:13
    .p1_wr_en   (_T_895),	// matmul/matmul-hw.mlir:17423:13
    .p1_wr_data (_T_894),	// matmul/matmul-hw.mlir:17424:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2356)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3280 (	// matmul/matmul-hw.mlir:17067:37
    .p0_rd_en   (_T_886),	// matmul/matmul-hw.mlir:17466:13
    .p1_wr_en   (_T_890),	// matmul/matmul-hw.mlir:17453:13
    .p1_wr_data (_T_889),	// matmul/matmul-hw.mlir:17454:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2355)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3281 (	// matmul/matmul-hw.mlir:17068:37
    .p0_rd_en   (_T_881),	// matmul/matmul-hw.mlir:17496:13
    .p1_wr_en   (_T_885),	// matmul/matmul-hw.mlir:17483:13
    .p1_wr_data (_T_884),	// matmul/matmul-hw.mlir:17484:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2354)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3282 (	// matmul/matmul-hw.mlir:17069:37
    .p0_rd_en   (_T_876),	// matmul/matmul-hw.mlir:17526:13
    .p1_wr_en   (_T_880),	// matmul/matmul-hw.mlir:17513:13
    .p1_wr_data (_T_879),	// matmul/matmul-hw.mlir:17514:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2353)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3283 (	// matmul/matmul-hw.mlir:17070:37
    .p0_rd_en   (_T_873),	// matmul/matmul-hw.mlir:17553:13
    .p1_wr_en   (_T_875),	// matmul/matmul-hw.mlir:17543:13
    .p1_wr_data (_T_874),	// matmul/matmul-hw.mlir:17544:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2352)
  );
  assign _T_955 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17071:13
  assign _T_954 = _T_2797 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8989:19, :17072:13
  assign _T_953 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17073:13
  assign _T_952 = _T_2786 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17074:13
  mult mult_inst80 (	// matmul/matmul-hw.mlir:17075:27
    .a      (A_reg_bank80_p0_rd_data),	// matmul/matmul-hw.mlir:12295:32
    .b      (_T_2459),
    .t      (_T_2786),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst80_result)
  );
  assign _T_951 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17076:13
  assign a_i_k_0_i_j_5 = A_reg_bank80_p0_rd_data;	// matmul/matmul-hw.mlir:12295:32, :17078:5
  //PROBE: a_i_k_0_i_j_5	// matmul/matmul-hw.mlir:17079:5
  assign b_i_k_0_i_j_5 = _T_2459;	// matmul/matmul-hw.mlir:17081:5
  //PROBE: b_i_k_0_i_j_5	// matmul/matmul-hw.mlir:17082:5
  assign c_prev_i_k_0_i_j_5 = C_reg_bank0_p0_rd_data_2368;	// matmul/matmul-hw.mlir:17054:36, :17084:5
  //PROBE: c_prev_i_k_0_i_j_5	// matmul/matmul-hw.mlir:17085:5
  assign tk_i_k_0_i_j_5 = _T_2764;	// matmul/matmul-hw.mlir:17087:5
  //PROBE: tk_i_k_0_i_j_5	// matmul/matmul-hw.mlir:17088:5
  wire [31:0] _T_3284 = mult_inst80_result + C_reg_bank0_p0_rd_data_2368;	// matmul/matmul-hw.mlir:17054:36, :17075:27, :17089:13
  assign c_i_k_0_i_j_5 = _T_3284;	// matmul/matmul-hw.mlir:17091:5
  //PROBE: c_i_k_0_i_j_5	// matmul/matmul-hw.mlir:17092:5
  assign _T_950 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17093:13
  assign _T_949 = _T_2808 ? _T_3284 : 32'bx;	// matmul/matmul-hw.mlir:8984:19, :17094:13
  localparam [3:0] _T_3286 = 4'h0;	// matmul/matmul-hw.mlir:17097:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17098:5
    if (rst)	// matmul/matmul-hw.mlir:17098:5
      i_k_next_3285 <= _T_3286;	// matmul/matmul-hw.mlir:17101:7
    else	// matmul/matmul-hw.mlir:17098:5
      i_k_next_3285 <= i_j_next_3265;	// matmul/matmul-hw.mlir:16979:13, :17099:7
  end // always @(posedge)
  assign _T_948 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17103:13
  assign _T_947 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17104:13
  mult mult_inst81 (	// matmul/matmul-hw.mlir:17105:27
    .a      (A_reg_bank81_p0_rd_data),	// matmul/matmul-hw.mlir:12296:32
    .b      (_T_2475),
    .t      (_T_2797),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst81_result)
  );
  assign _T_946 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17106:13
  assign a_i_k_1_i_j_5 = A_reg_bank81_p0_rd_data;	// matmul/matmul-hw.mlir:12296:32, :17108:5
  //PROBE: a_i_k_1_i_j_5	// matmul/matmul-hw.mlir:17109:5
  assign b_i_k_1_i_j_5 = _T_2475;	// matmul/matmul-hw.mlir:17111:5
  //PROBE: b_i_k_1_i_j_5	// matmul/matmul-hw.mlir:17112:5
  assign c_prev_i_k_1_i_j_5 = C_reg_bank1_p0_rd_data_2367;	// matmul/matmul-hw.mlir:17055:36, :17114:5
  //PROBE: c_prev_i_k_1_i_j_5	// matmul/matmul-hw.mlir:17115:5
  assign tk_i_k_1_i_j_5 = _T_2775;	// matmul/matmul-hw.mlir:17117:5
  //PROBE: tk_i_k_1_i_j_5	// matmul/matmul-hw.mlir:17118:5
  wire [31:0] _T_3287 = mult_inst81_result + C_reg_bank1_p0_rd_data_2367;	// matmul/matmul-hw.mlir:17055:36, :17105:27, :17119:13
  assign c_i_k_1_i_j_5 = _T_3287;	// matmul/matmul-hw.mlir:17121:5
  //PROBE: c_i_k_1_i_j_5	// matmul/matmul-hw.mlir:17122:5
  assign _T_945 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17123:13
  assign _T_944 = _T_2819 ? _T_3287 : 32'bx;	// matmul/matmul-hw.mlir:8979:19, :17124:13
  localparam [3:0] _T_3289 = 4'h0;	// matmul/matmul-hw.mlir:17127:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17128:5
    if (rst)	// matmul/matmul-hw.mlir:17128:5
      i_k_next_3288 <= _T_3289;	// matmul/matmul-hw.mlir:17131:7
    else	// matmul/matmul-hw.mlir:17128:5
      i_k_next_3288 <= i_k_next_3285;	// matmul/matmul-hw.mlir:17096:13, :17129:7
  end // always @(posedge)
  assign _T_943 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17133:13
  assign _T_942 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17134:13
  mult mult_inst82 (	// matmul/matmul-hw.mlir:17135:27
    .a      (A_reg_bank82_p0_rd_data),	// matmul/matmul-hw.mlir:12297:32
    .b      (_T_2491),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst82_result)
  );
  assign _T_941 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17136:13
  assign a_i_k_2_i_j_5 = A_reg_bank82_p0_rd_data;	// matmul/matmul-hw.mlir:12297:32, :17138:5
  //PROBE: a_i_k_2_i_j_5	// matmul/matmul-hw.mlir:17139:5
  assign b_i_k_2_i_j_5 = _T_2491;	// matmul/matmul-hw.mlir:17141:5
  //PROBE: b_i_k_2_i_j_5	// matmul/matmul-hw.mlir:17142:5
  assign c_prev_i_k_2_i_j_5 = C_reg_bank2_p0_rd_data_2366;	// matmul/matmul-hw.mlir:17056:36, :17144:5
  //PROBE: c_prev_i_k_2_i_j_5	// matmul/matmul-hw.mlir:17145:5
  assign tk_i_k_2_i_j_5 = _T_2786;	// matmul/matmul-hw.mlir:17147:5
  //PROBE: tk_i_k_2_i_j_5	// matmul/matmul-hw.mlir:17148:5
  wire [31:0] _T_3290 = mult_inst82_result + C_reg_bank2_p0_rd_data_2366;	// matmul/matmul-hw.mlir:17056:36, :17135:27, :17149:13
  assign c_i_k_2_i_j_5 = _T_3290;	// matmul/matmul-hw.mlir:17151:5
  //PROBE: c_i_k_2_i_j_5	// matmul/matmul-hw.mlir:17152:5
  assign _T_940 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17153:13
  assign _T_939 = _T_2830 ? _T_3290 : 32'bx;	// matmul/matmul-hw.mlir:8974:19, :17154:13
  localparam [3:0] _T_3292 = 4'h0;	// matmul/matmul-hw.mlir:17157:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17158:5
    if (rst)	// matmul/matmul-hw.mlir:17158:5
      i_k_next_3291 <= _T_3292;	// matmul/matmul-hw.mlir:17161:7
    else	// matmul/matmul-hw.mlir:17158:5
      i_k_next_3291 <= i_k_next_3288;	// matmul/matmul-hw.mlir:17126:13, :17159:7
  end // always @(posedge)
  assign _T_938 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17163:13
  assign _T_937 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17164:13
  mult mult_inst83 (	// matmul/matmul-hw.mlir:17165:27
    .a      (A_reg_bank83_p0_rd_data),	// matmul/matmul-hw.mlir:12298:32
    .b      (_T_2507),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst83_result)
  );
  assign _T_936 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17166:13
  assign a_i_k_3_i_j_5 = A_reg_bank83_p0_rd_data;	// matmul/matmul-hw.mlir:12298:32, :17168:5
  //PROBE: a_i_k_3_i_j_5	// matmul/matmul-hw.mlir:17169:5
  assign b_i_k_3_i_j_5 = _T_2507;	// matmul/matmul-hw.mlir:17171:5
  //PROBE: b_i_k_3_i_j_5	// matmul/matmul-hw.mlir:17172:5
  assign c_prev_i_k_3_i_j_5 = C_reg_bank3_p0_rd_data_2365;	// matmul/matmul-hw.mlir:17057:36, :17174:5
  //PROBE: c_prev_i_k_3_i_j_5	// matmul/matmul-hw.mlir:17175:5
  assign tk_i_k_3_i_j_5 = _T_2797;	// matmul/matmul-hw.mlir:17177:5
  //PROBE: tk_i_k_3_i_j_5	// matmul/matmul-hw.mlir:17178:5
  wire [31:0] _T_3293 = mult_inst83_result + C_reg_bank3_p0_rd_data_2365;	// matmul/matmul-hw.mlir:17057:36, :17165:27, :17179:13
  assign c_i_k_3_i_j_5 = _T_3293;	// matmul/matmul-hw.mlir:17181:5
  //PROBE: c_i_k_3_i_j_5	// matmul/matmul-hw.mlir:17182:5
  assign _T_935 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17183:13
  assign _T_934 = _T_2841 ? _T_3293 : 32'bx;	// matmul/matmul-hw.mlir:8969:19, :17184:13
  localparam [3:0] _T_3295 = 4'h0;	// matmul/matmul-hw.mlir:17187:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17188:5
    if (rst)	// matmul/matmul-hw.mlir:17188:5
      i_k_next_3294 <= _T_3295;	// matmul/matmul-hw.mlir:17191:7
    else	// matmul/matmul-hw.mlir:17188:5
      i_k_next_3294 <= i_k_next_3291;	// matmul/matmul-hw.mlir:17156:13, :17189:7
  end // always @(posedge)
  assign _T_933 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17193:13
  assign _T_932 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17194:13
  mult mult_inst84 (	// matmul/matmul-hw.mlir:17195:27
    .a      (A_reg_bank84_p0_rd_data),	// matmul/matmul-hw.mlir:12299:32
    .b      (_T_2523),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst84_result)
  );
  assign _T_931 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17196:13
  assign a_i_k_4_i_j_5 = A_reg_bank84_p0_rd_data;	// matmul/matmul-hw.mlir:12299:32, :17198:5
  //PROBE: a_i_k_4_i_j_5	// matmul/matmul-hw.mlir:17199:5
  assign b_i_k_4_i_j_5 = _T_2523;	// matmul/matmul-hw.mlir:17201:5
  //PROBE: b_i_k_4_i_j_5	// matmul/matmul-hw.mlir:17202:5
  assign c_prev_i_k_4_i_j_5 = C_reg_bank4_p0_rd_data_2364;	// matmul/matmul-hw.mlir:17058:36, :17204:5
  //PROBE: c_prev_i_k_4_i_j_5	// matmul/matmul-hw.mlir:17205:5
  assign tk_i_k_4_i_j_5 = _T_2808;	// matmul/matmul-hw.mlir:17207:5
  //PROBE: tk_i_k_4_i_j_5	// matmul/matmul-hw.mlir:17208:5
  wire [31:0] _T_3296 = mult_inst84_result + C_reg_bank4_p0_rd_data_2364;	// matmul/matmul-hw.mlir:17058:36, :17195:27, :17209:13
  assign c_i_k_4_i_j_5 = _T_3296;	// matmul/matmul-hw.mlir:17211:5
  //PROBE: c_i_k_4_i_j_5	// matmul/matmul-hw.mlir:17212:5
  assign _T_930 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17213:13
  assign _T_929 = _T_2852 ? _T_3296 : 32'bx;	// matmul/matmul-hw.mlir:8964:19, :17214:13
  localparam [3:0] _T_3298 = 4'h0;	// matmul/matmul-hw.mlir:17217:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17218:5
    if (rst)	// matmul/matmul-hw.mlir:17218:5
      i_k_next_3297 <= _T_3298;	// matmul/matmul-hw.mlir:17221:7
    else	// matmul/matmul-hw.mlir:17218:5
      i_k_next_3297 <= i_k_next_3294;	// matmul/matmul-hw.mlir:17186:13, :17219:7
  end // always @(posedge)
  assign _T_928 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17223:13
  assign _T_927 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17224:13
  mult mult_inst85 (	// matmul/matmul-hw.mlir:17225:27
    .a      (A_reg_bank85_p0_rd_data),	// matmul/matmul-hw.mlir:12300:32
    .b      (_T_2539),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst85_result)
  );
  assign _T_926 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17226:13
  assign a_i_k_5_i_j_5 = A_reg_bank85_p0_rd_data;	// matmul/matmul-hw.mlir:12300:32, :17228:5
  //PROBE: a_i_k_5_i_j_5	// matmul/matmul-hw.mlir:17229:5
  assign b_i_k_5_i_j_5 = _T_2539;	// matmul/matmul-hw.mlir:17231:5
  //PROBE: b_i_k_5_i_j_5	// matmul/matmul-hw.mlir:17232:5
  assign c_prev_i_k_5_i_j_5 = C_reg_bank5_p0_rd_data_2363;	// matmul/matmul-hw.mlir:17059:36, :17234:5
  //PROBE: c_prev_i_k_5_i_j_5	// matmul/matmul-hw.mlir:17235:5
  assign tk_i_k_5_i_j_5 = _T_2819;	// matmul/matmul-hw.mlir:17237:5
  //PROBE: tk_i_k_5_i_j_5	// matmul/matmul-hw.mlir:17238:5
  wire [31:0] _T_3299 = mult_inst85_result + C_reg_bank5_p0_rd_data_2363;	// matmul/matmul-hw.mlir:17059:36, :17225:27, :17239:13
  assign c_i_k_5_i_j_5 = _T_3299;	// matmul/matmul-hw.mlir:17241:5
  //PROBE: c_i_k_5_i_j_5	// matmul/matmul-hw.mlir:17242:5
  assign _T_925 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17243:13
  assign _T_924 = _T_2863 ? _T_3299 : 32'bx;	// matmul/matmul-hw.mlir:8959:19, :17244:13
  localparam [3:0] _T_3301 = 4'h0;	// matmul/matmul-hw.mlir:17247:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17248:5
    if (rst)	// matmul/matmul-hw.mlir:17248:5
      i_k_next_3300 <= _T_3301;	// matmul/matmul-hw.mlir:17251:7
    else	// matmul/matmul-hw.mlir:17248:5
      i_k_next_3300 <= i_k_next_3297;	// matmul/matmul-hw.mlir:17216:13, :17249:7
  end // always @(posedge)
  assign _T_923 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17253:13
  assign _T_922 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17254:13
  mult mult_inst86 (	// matmul/matmul-hw.mlir:17255:27
    .a      (A_reg_bank86_p0_rd_data),	// matmul/matmul-hw.mlir:12301:32
    .b      (_T_2555),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst86_result)
  );
  assign _T_921 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17256:13
  assign a_i_k_6_i_j_5 = A_reg_bank86_p0_rd_data;	// matmul/matmul-hw.mlir:12301:32, :17258:5
  //PROBE: a_i_k_6_i_j_5	// matmul/matmul-hw.mlir:17259:5
  assign b_i_k_6_i_j_5 = _T_2555;	// matmul/matmul-hw.mlir:17261:5
  //PROBE: b_i_k_6_i_j_5	// matmul/matmul-hw.mlir:17262:5
  assign c_prev_i_k_6_i_j_5 = C_reg_bank6_p0_rd_data_2362;	// matmul/matmul-hw.mlir:17060:36, :17264:5
  //PROBE: c_prev_i_k_6_i_j_5	// matmul/matmul-hw.mlir:17265:5
  assign tk_i_k_6_i_j_5 = _T_2830;	// matmul/matmul-hw.mlir:17267:5
  //PROBE: tk_i_k_6_i_j_5	// matmul/matmul-hw.mlir:17268:5
  wire [31:0] _T_3302 = mult_inst86_result + C_reg_bank6_p0_rd_data_2362;	// matmul/matmul-hw.mlir:17060:36, :17255:27, :17269:13
  assign c_i_k_6_i_j_5 = _T_3302;	// matmul/matmul-hw.mlir:17271:5
  //PROBE: c_i_k_6_i_j_5	// matmul/matmul-hw.mlir:17272:5
  assign _T_920 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17273:13
  assign _T_919 = _T_2874 ? _T_3302 : 32'bx;	// matmul/matmul-hw.mlir:8954:19, :17274:13
  localparam [3:0] _T_3304 = 4'h0;	// matmul/matmul-hw.mlir:17277:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17278:5
    if (rst)	// matmul/matmul-hw.mlir:17278:5
      i_k_next_3303 <= _T_3304;	// matmul/matmul-hw.mlir:17281:7
    else	// matmul/matmul-hw.mlir:17278:5
      i_k_next_3303 <= i_k_next_3300;	// matmul/matmul-hw.mlir:17246:13, :17279:7
  end // always @(posedge)
  assign _T_918 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17283:13
  assign _T_917 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17284:13
  mult mult_inst87 (	// matmul/matmul-hw.mlir:17285:27
    .a      (A_reg_bank87_p0_rd_data),	// matmul/matmul-hw.mlir:12302:32
    .b      (_T_2571),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst87_result)
  );
  assign _T_916 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17286:13
  assign a_i_k_7_i_j_5 = A_reg_bank87_p0_rd_data;	// matmul/matmul-hw.mlir:12302:32, :17288:5
  //PROBE: a_i_k_7_i_j_5	// matmul/matmul-hw.mlir:17289:5
  assign b_i_k_7_i_j_5 = _T_2571;	// matmul/matmul-hw.mlir:17291:5
  //PROBE: b_i_k_7_i_j_5	// matmul/matmul-hw.mlir:17292:5
  assign c_prev_i_k_7_i_j_5 = C_reg_bank7_p0_rd_data_2361;	// matmul/matmul-hw.mlir:17061:36, :17294:5
  //PROBE: c_prev_i_k_7_i_j_5	// matmul/matmul-hw.mlir:17295:5
  assign tk_i_k_7_i_j_5 = _T_2841;	// matmul/matmul-hw.mlir:17297:5
  //PROBE: tk_i_k_7_i_j_5	// matmul/matmul-hw.mlir:17298:5
  wire [31:0] _T_3305 = mult_inst87_result + C_reg_bank7_p0_rd_data_2361;	// matmul/matmul-hw.mlir:17061:36, :17285:27, :17299:13
  assign c_i_k_7_i_j_5 = _T_3305;	// matmul/matmul-hw.mlir:17301:5
  //PROBE: c_i_k_7_i_j_5	// matmul/matmul-hw.mlir:17302:5
  assign _T_915 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17303:13
  assign _T_914 = _T_2885 ? _T_3305 : 32'bx;	// matmul/matmul-hw.mlir:8949:19, :17304:13
  localparam [3:0] _T_3307 = 4'h0;	// matmul/matmul-hw.mlir:17307:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17308:5
    if (rst)	// matmul/matmul-hw.mlir:17308:5
      i_k_next_3306 <= _T_3307;	// matmul/matmul-hw.mlir:17311:7
    else	// matmul/matmul-hw.mlir:17308:5
      i_k_next_3306 <= i_k_next_3303;	// matmul/matmul-hw.mlir:17276:13, :17309:7
  end // always @(posedge)
  assign _T_913 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17313:13
  assign _T_912 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17314:13
  mult mult_inst88 (	// matmul/matmul-hw.mlir:17315:27
    .a      (A_reg_bank88_p0_rd_data),	// matmul/matmul-hw.mlir:12303:32
    .b      (_T_2587),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst88_result)
  );
  assign _T_911 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17316:13
  assign a_i_k_8_i_j_5 = A_reg_bank88_p0_rd_data;	// matmul/matmul-hw.mlir:12303:32, :17318:5
  //PROBE: a_i_k_8_i_j_5	// matmul/matmul-hw.mlir:17319:5
  assign b_i_k_8_i_j_5 = _T_2587;	// matmul/matmul-hw.mlir:17321:5
  //PROBE: b_i_k_8_i_j_5	// matmul/matmul-hw.mlir:17322:5
  assign c_prev_i_k_8_i_j_5 = C_reg_bank8_p0_rd_data_2360;	// matmul/matmul-hw.mlir:17062:36, :17324:5
  //PROBE: c_prev_i_k_8_i_j_5	// matmul/matmul-hw.mlir:17325:5
  assign tk_i_k_8_i_j_5 = _T_2852;	// matmul/matmul-hw.mlir:17327:5
  //PROBE: tk_i_k_8_i_j_5	// matmul/matmul-hw.mlir:17328:5
  wire [31:0] _T_3308 = mult_inst88_result + C_reg_bank8_p0_rd_data_2360;	// matmul/matmul-hw.mlir:17062:36, :17315:27, :17329:13
  assign c_i_k_8_i_j_5 = _T_3308;	// matmul/matmul-hw.mlir:17331:5
  //PROBE: c_i_k_8_i_j_5	// matmul/matmul-hw.mlir:17332:5
  assign _T_910 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17333:13
  assign _T_909 = _T_2892 ? _T_3308 : 32'bx;	// matmul/matmul-hw.mlir:8944:19, :17334:13
  localparam [3:0] _T_3310 = 4'h0;	// matmul/matmul-hw.mlir:17337:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17338:5
    if (rst)	// matmul/matmul-hw.mlir:17338:5
      i_k_next_3309 <= _T_3310;	// matmul/matmul-hw.mlir:17341:7
    else	// matmul/matmul-hw.mlir:17338:5
      i_k_next_3309 <= i_k_next_3306;	// matmul/matmul-hw.mlir:17306:13, :17339:7
  end // always @(posedge)
  assign _T_908 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17343:13
  assign _T_907 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17344:13
  mult mult_inst89 (	// matmul/matmul-hw.mlir:17345:27
    .a      (A_reg_bank89_p0_rd_data),	// matmul/matmul-hw.mlir:12304:32
    .b      (_T_2603),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst89_result)
  );
  assign _T_906 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17346:13
  assign a_i_k_9_i_j_5 = A_reg_bank89_p0_rd_data;	// matmul/matmul-hw.mlir:12304:32, :17348:5
  //PROBE: a_i_k_9_i_j_5	// matmul/matmul-hw.mlir:17349:5
  assign b_i_k_9_i_j_5 = _T_2603;	// matmul/matmul-hw.mlir:17351:5
  //PROBE: b_i_k_9_i_j_5	// matmul/matmul-hw.mlir:17352:5
  assign c_prev_i_k_9_i_j_5 = C_reg_bank9_p0_rd_data_2359;	// matmul/matmul-hw.mlir:17063:36, :17354:5
  //PROBE: c_prev_i_k_9_i_j_5	// matmul/matmul-hw.mlir:17355:5
  assign tk_i_k_9_i_j_5 = _T_2863;	// matmul/matmul-hw.mlir:17357:5
  //PROBE: tk_i_k_9_i_j_5	// matmul/matmul-hw.mlir:17358:5
  wire [31:0] _T_3311 = mult_inst89_result + C_reg_bank9_p0_rd_data_2359;	// matmul/matmul-hw.mlir:17063:36, :17345:27, :17359:13
  assign c_i_k_9_i_j_5 = _T_3311;	// matmul/matmul-hw.mlir:17361:5
  //PROBE: c_i_k_9_i_j_5	// matmul/matmul-hw.mlir:17362:5
  assign _T_905 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17363:13
  assign _T_904 = _T_2897 ? _T_3311 : 32'bx;	// matmul/matmul-hw.mlir:8939:19, :17364:13
  localparam [3:0] _T_3313 = 4'h0;	// matmul/matmul-hw.mlir:17367:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17368:5
    if (rst)	// matmul/matmul-hw.mlir:17368:5
      i_k_next_3312 <= _T_3313;	// matmul/matmul-hw.mlir:17371:7
    else	// matmul/matmul-hw.mlir:17368:5
      i_k_next_3312 <= i_k_next_3309;	// matmul/matmul-hw.mlir:17336:13, :17369:7
  end // always @(posedge)
  assign _T_903 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17373:13
  assign _T_902 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17374:13
  mult mult_inst90 (	// matmul/matmul-hw.mlir:17375:27
    .a      (A_reg_bank90_p0_rd_data),	// matmul/matmul-hw.mlir:12305:32
    .b      (_T_2619),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst90_result)
  );
  assign _T_901 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17376:13
  assign a_i_k_10_i_j_5 = A_reg_bank90_p0_rd_data;	// matmul/matmul-hw.mlir:12305:32, :17378:5
  //PROBE: a_i_k_10_i_j_5	// matmul/matmul-hw.mlir:17379:5
  assign b_i_k_10_i_j_5 = _T_2619;	// matmul/matmul-hw.mlir:17381:5
  //PROBE: b_i_k_10_i_j_5	// matmul/matmul-hw.mlir:17382:5
  assign c_prev_i_k_10_i_j_5 = C_reg_bank10_p0_rd_data_2358;	// matmul/matmul-hw.mlir:17064:37, :17384:5
  //PROBE: c_prev_i_k_10_i_j_5	// matmul/matmul-hw.mlir:17385:5
  assign tk_i_k_10_i_j_5 = _T_2874;	// matmul/matmul-hw.mlir:17387:5
  //PROBE: tk_i_k_10_i_j_5	// matmul/matmul-hw.mlir:17388:5
  wire [31:0] _T_3314 = mult_inst90_result + C_reg_bank10_p0_rd_data_2358;	// matmul/matmul-hw.mlir:17064:37, :17375:27, :17389:13
  assign c_i_k_10_i_j_5 = _T_3314;	// matmul/matmul-hw.mlir:17391:5
  //PROBE: c_i_k_10_i_j_5	// matmul/matmul-hw.mlir:17392:5
  assign _T_900 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17393:13
  assign _T_899 = _T_2902 ? _T_3314 : 32'bx;	// matmul/matmul-hw.mlir:8934:19, :17394:13
  localparam [3:0] _T_3316 = 4'h0;	// matmul/matmul-hw.mlir:17397:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17398:5
    if (rst)	// matmul/matmul-hw.mlir:17398:5
      i_k_next_3315 <= _T_3316;	// matmul/matmul-hw.mlir:17401:7
    else	// matmul/matmul-hw.mlir:17398:5
      i_k_next_3315 <= i_k_next_3312;	// matmul/matmul-hw.mlir:17366:13, :17399:7
  end // always @(posedge)
  assign _T_898 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17403:13
  assign _T_897 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17404:13
  mult mult_inst91 (	// matmul/matmul-hw.mlir:17405:27
    .a      (A_reg_bank91_p0_rd_data),	// matmul/matmul-hw.mlir:12306:32
    .b      (_T_2635),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst91_result)
  );
  assign _T_896 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17406:13
  assign a_i_k_11_i_j_5 = A_reg_bank91_p0_rd_data;	// matmul/matmul-hw.mlir:12306:32, :17408:5
  //PROBE: a_i_k_11_i_j_5	// matmul/matmul-hw.mlir:17409:5
  assign b_i_k_11_i_j_5 = _T_2635;	// matmul/matmul-hw.mlir:17411:5
  //PROBE: b_i_k_11_i_j_5	// matmul/matmul-hw.mlir:17412:5
  assign c_prev_i_k_11_i_j_5 = C_reg_bank11_p0_rd_data_2357;	// matmul/matmul-hw.mlir:17065:37, :17414:5
  //PROBE: c_prev_i_k_11_i_j_5	// matmul/matmul-hw.mlir:17415:5
  assign tk_i_k_11_i_j_5 = _T_2885;	// matmul/matmul-hw.mlir:17417:5
  //PROBE: tk_i_k_11_i_j_5	// matmul/matmul-hw.mlir:17418:5
  wire [31:0] _T_3317 = mult_inst91_result + C_reg_bank11_p0_rd_data_2357;	// matmul/matmul-hw.mlir:17065:37, :17405:27, :17419:13
  assign c_i_k_11_i_j_5 = _T_3317;	// matmul/matmul-hw.mlir:17421:5
  //PROBE: c_i_k_11_i_j_5	// matmul/matmul-hw.mlir:17422:5
  assign _T_895 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17423:13
  assign _T_894 = _T_2907 ? _T_3317 : 32'bx;	// matmul/matmul-hw.mlir:8929:19, :17424:13
  localparam [3:0] _T_3319 = 4'h0;	// matmul/matmul-hw.mlir:17427:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17428:5
    if (rst)	// matmul/matmul-hw.mlir:17428:5
      i_k_next_3318 <= _T_3319;	// matmul/matmul-hw.mlir:17431:7
    else	// matmul/matmul-hw.mlir:17428:5
      i_k_next_3318 <= i_k_next_3315;	// matmul/matmul-hw.mlir:17396:13, :17429:7
  end // always @(posedge)
  assign _T_893 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17433:13
  assign _T_892 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17434:13
  mult mult_inst92 (	// matmul/matmul-hw.mlir:17435:27
    .a      (A_reg_bank92_p0_rd_data),	// matmul/matmul-hw.mlir:12307:32
    .b      (_T_2651),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst92_result)
  );
  assign _T_891 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17436:13
  assign a_i_k_12_i_j_5 = A_reg_bank92_p0_rd_data;	// matmul/matmul-hw.mlir:12307:32, :17438:5
  //PROBE: a_i_k_12_i_j_5	// matmul/matmul-hw.mlir:17439:5
  assign b_i_k_12_i_j_5 = _T_2651;	// matmul/matmul-hw.mlir:17441:5
  //PROBE: b_i_k_12_i_j_5	// matmul/matmul-hw.mlir:17442:5
  assign c_prev_i_k_12_i_j_5 = C_reg_bank12_p0_rd_data_2356;	// matmul/matmul-hw.mlir:17066:37, :17444:5
  //PROBE: c_prev_i_k_12_i_j_5	// matmul/matmul-hw.mlir:17445:5
  assign tk_i_k_12_i_j_5 = _T_2892;	// matmul/matmul-hw.mlir:17447:5
  //PROBE: tk_i_k_12_i_j_5	// matmul/matmul-hw.mlir:17448:5
  wire [31:0] _T_3320 = mult_inst92_result + C_reg_bank12_p0_rd_data_2356;	// matmul/matmul-hw.mlir:17066:37, :17435:27, :17449:13
  assign c_i_k_12_i_j_5 = _T_3320;	// matmul/matmul-hw.mlir:17451:5
  //PROBE: c_i_k_12_i_j_5	// matmul/matmul-hw.mlir:17452:5
  assign _T_890 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17453:13
  assign _T_889 = _T_2912 ? _T_3320 : 32'bx;	// matmul/matmul-hw.mlir:8924:19, :17454:13
  localparam [3:0] _T_3322 = 4'h0;	// matmul/matmul-hw.mlir:17457:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17458:5
    if (rst)	// matmul/matmul-hw.mlir:17458:5
      i_k_next_3321 <= _T_3322;	// matmul/matmul-hw.mlir:17461:7
    else	// matmul/matmul-hw.mlir:17458:5
      i_k_next_3321 <= i_k_next_3318;	// matmul/matmul-hw.mlir:17426:13, :17459:7
  end // always @(posedge)
  assign _T_888 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17463:13
  assign _T_887 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17464:13
  mult mult_inst93 (	// matmul/matmul-hw.mlir:17465:27
    .a      (A_reg_bank93_p0_rd_data),	// matmul/matmul-hw.mlir:12308:32
    .b      (_T_2667),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst93_result)
  );
  assign _T_886 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17466:13
  assign a_i_k_13_i_j_5 = A_reg_bank93_p0_rd_data;	// matmul/matmul-hw.mlir:12308:32, :17468:5
  //PROBE: a_i_k_13_i_j_5	// matmul/matmul-hw.mlir:17469:5
  assign b_i_k_13_i_j_5 = _T_2667;	// matmul/matmul-hw.mlir:17471:5
  //PROBE: b_i_k_13_i_j_5	// matmul/matmul-hw.mlir:17472:5
  assign c_prev_i_k_13_i_j_5 = C_reg_bank13_p0_rd_data_2355;	// matmul/matmul-hw.mlir:17067:37, :17474:5
  //PROBE: c_prev_i_k_13_i_j_5	// matmul/matmul-hw.mlir:17475:5
  assign tk_i_k_13_i_j_5 = _T_2897;	// matmul/matmul-hw.mlir:17477:5
  //PROBE: tk_i_k_13_i_j_5	// matmul/matmul-hw.mlir:17478:5
  wire [31:0] _T_3323 = mult_inst93_result + C_reg_bank13_p0_rd_data_2355;	// matmul/matmul-hw.mlir:17067:37, :17465:27, :17479:13
  assign c_i_k_13_i_j_5 = _T_3323;	// matmul/matmul-hw.mlir:17481:5
  //PROBE: c_i_k_13_i_j_5	// matmul/matmul-hw.mlir:17482:5
  assign _T_885 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17483:13
  assign _T_884 = _T_2917 ? _T_3323 : 32'bx;	// matmul/matmul-hw.mlir:8919:19, :17484:13
  localparam [3:0] _T_3325 = 4'h0;	// matmul/matmul-hw.mlir:17487:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17488:5
    if (rst)	// matmul/matmul-hw.mlir:17488:5
      i_k_next_3324 <= _T_3325;	// matmul/matmul-hw.mlir:17491:7
    else	// matmul/matmul-hw.mlir:17488:5
      i_k_next_3324 <= i_k_next_3321;	// matmul/matmul-hw.mlir:17456:13, :17489:7
  end // always @(posedge)
  assign _T_883 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17493:13
  assign _T_882 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17494:13
  mult mult_inst94 (	// matmul/matmul-hw.mlir:17495:27
    .a      (A_reg_bank94_p0_rd_data),	// matmul/matmul-hw.mlir:12309:32
    .b      (_T_2683),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst94_result)
  );
  assign _T_881 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17496:13
  assign a_i_k_14_i_j_5 = A_reg_bank94_p0_rd_data;	// matmul/matmul-hw.mlir:12309:32, :17498:5
  //PROBE: a_i_k_14_i_j_5	// matmul/matmul-hw.mlir:17499:5
  assign b_i_k_14_i_j_5 = _T_2683;	// matmul/matmul-hw.mlir:17501:5
  //PROBE: b_i_k_14_i_j_5	// matmul/matmul-hw.mlir:17502:5
  assign c_prev_i_k_14_i_j_5 = C_reg_bank14_p0_rd_data_2354;	// matmul/matmul-hw.mlir:17068:37, :17504:5
  //PROBE: c_prev_i_k_14_i_j_5	// matmul/matmul-hw.mlir:17505:5
  assign tk_i_k_14_i_j_5 = _T_2902;	// matmul/matmul-hw.mlir:17507:5
  //PROBE: tk_i_k_14_i_j_5	// matmul/matmul-hw.mlir:17508:5
  wire [31:0] _T_3326 = mult_inst94_result + C_reg_bank14_p0_rd_data_2354;	// matmul/matmul-hw.mlir:17068:37, :17495:27, :17509:13
  assign c_i_k_14_i_j_5 = _T_3326;	// matmul/matmul-hw.mlir:17511:5
  //PROBE: c_i_k_14_i_j_5	// matmul/matmul-hw.mlir:17512:5
  assign _T_880 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17513:13
  assign _T_879 = _T_2922 ? _T_3326 : 32'bx;	// matmul/matmul-hw.mlir:8914:19, :17514:13
  localparam [3:0] _T_3328 = 4'h0;	// matmul/matmul-hw.mlir:17517:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17518:5
    if (rst)	// matmul/matmul-hw.mlir:17518:5
      i_k_next_3327 <= _T_3328;	// matmul/matmul-hw.mlir:17521:7
    else	// matmul/matmul-hw.mlir:17518:5
      i_k_next_3327 <= i_k_next_3324;	// matmul/matmul-hw.mlir:17486:13, :17519:7
  end // always @(posedge)
  assign _T_878 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17523:13
  assign _T_877 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17524:13
  mult mult_inst95 (	// matmul/matmul-hw.mlir:17525:27
    .a      (A_reg_bank95_p0_rd_data),	// matmul/matmul-hw.mlir:12310:32
    .b      (_T_2699),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst95_result)
  );
  assign _T_876 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17526:13
  assign a_i_k_15_i_j_5 = A_reg_bank95_p0_rd_data;	// matmul/matmul-hw.mlir:12310:32, :17528:5
  //PROBE: a_i_k_15_i_j_5	// matmul/matmul-hw.mlir:17529:5
  assign b_i_k_15_i_j_5 = _T_2699;	// matmul/matmul-hw.mlir:17531:5
  //PROBE: b_i_k_15_i_j_5	// matmul/matmul-hw.mlir:17532:5
  assign c_prev_i_k_15_i_j_5 = C_reg_bank15_p0_rd_data_2353;	// matmul/matmul-hw.mlir:17069:37, :17534:5
  //PROBE: c_prev_i_k_15_i_j_5	// matmul/matmul-hw.mlir:17535:5
  assign tk_i_k_15_i_j_5 = _T_2907;	// matmul/matmul-hw.mlir:17537:5
  //PROBE: tk_i_k_15_i_j_5	// matmul/matmul-hw.mlir:17538:5
  wire [31:0] _T_3329 = mult_inst95_result + C_reg_bank15_p0_rd_data_2353;	// matmul/matmul-hw.mlir:17069:37, :17525:27, :17539:13
  assign c_i_k_15_i_j_5 = _T_3329;	// matmul/matmul-hw.mlir:17541:5
  //PROBE: c_i_k_15_i_j_5	// matmul/matmul-hw.mlir:17542:5
  assign _T_875 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17543:13
  assign _T_874 = _T_2927 ? _T_3329 : 32'bx;	// matmul/matmul-hw.mlir:8909:19, :17544:13
  localparam [3:0] _T_3331 = 4'h0;	// matmul/matmul-hw.mlir:17547:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17548:5
    if (rst)	// matmul/matmul-hw.mlir:17548:5
      i_k_next_3330 <= _T_3331;	// matmul/matmul-hw.mlir:17551:7
    else	// matmul/matmul-hw.mlir:17548:5
      i_k_next_3330 <= i_k_next_3327;	// matmul/matmul-hw.mlir:17516:13, :17549:7
  end // always @(posedge)
  assign _T_873 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17553:13
  wire [3:0][3:0] _T_3333 = i_delayed_3332;	// matmul/matmul-hw.mlir:17555:13
  wire [3:0][3:0] _T_3334 = {_T_3333[2'h0+:3], {{i_k_next_3330}}};	// matmul/matmul-hw.mlir:17546:13, :17556:19, :17557:13, :17558:13, :17559:13
  wire [3:0][3:0] _T_3335 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:17560:19, :17561:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17562:5
    if (rst)	// matmul/matmul-hw.mlir:17562:5
      i_delayed_3332 <= _T_3335;	// matmul/matmul-hw.mlir:17565:7
    else	// matmul/matmul-hw.mlir:17562:5
      i_delayed_3332 <= _T_3334;	// matmul/matmul-hw.mlir:17563:7
  end // always @(posedge)
  assign _T_872 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17569:13
  assign _T_871 = _T_2932 ? i_delayed_3332[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8906:18, :17555:13, :17567:20, :17568:13, :17570:13
  assign _T_870 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17571:13
  assign _T_869 = _T_2932 ? C_reg_bank16_p0_rd_data_2352 : 32'bx;	// matmul/matmul-hw.mlir:8904:19, :17070:37, :17572:13
  localparam [3:0] _T_3337 = 4'h0;	// matmul/matmul-hw.mlir:17575:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17576:5
    if (rst)	// matmul/matmul-hw.mlir:17576:5
      i_j_next_3336 <= _T_3337;	// matmul/matmul-hw.mlir:17579:7
    else	// matmul/matmul-hw.mlir:17576:5
      i_j_next_3336 <= i_j_next_3265;	// matmul/matmul-hw.mlir:16979:13, :17577:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3338 (	// matmul/matmul-hw.mlir:17649:36
    .p0_rd_en   (_T_864),	// matmul/matmul-hw.mlir:17671:13
    .p1_wr_en   (_T_868),	// matmul/matmul-hw.mlir:17666:13
    .p1_wr_data (_T_867),	// matmul/matmul-hw.mlir:17667:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2351)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3339 (	// matmul/matmul-hw.mlir:17650:36
    .p0_rd_en   (_T_859),	// matmul/matmul-hw.mlir:17701:13
    .p1_wr_en   (_T_863),	// matmul/matmul-hw.mlir:17688:13
    .p1_wr_data (_T_862),	// matmul/matmul-hw.mlir:17689:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2350)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3340 (	// matmul/matmul-hw.mlir:17651:36
    .p0_rd_en   (_T_854),	// matmul/matmul-hw.mlir:17731:13
    .p1_wr_en   (_T_858),	// matmul/matmul-hw.mlir:17718:13
    .p1_wr_data (_T_857),	// matmul/matmul-hw.mlir:17719:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2349)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3341 (	// matmul/matmul-hw.mlir:17652:36
    .p0_rd_en   (_T_849),	// matmul/matmul-hw.mlir:17761:13
    .p1_wr_en   (_T_853),	// matmul/matmul-hw.mlir:17748:13
    .p1_wr_data (_T_852),	// matmul/matmul-hw.mlir:17749:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2348)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3342 (	// matmul/matmul-hw.mlir:17653:36
    .p0_rd_en   (_T_844),	// matmul/matmul-hw.mlir:17791:13
    .p1_wr_en   (_T_848),	// matmul/matmul-hw.mlir:17778:13
    .p1_wr_data (_T_847),	// matmul/matmul-hw.mlir:17779:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2347)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3343 (	// matmul/matmul-hw.mlir:17654:36
    .p0_rd_en   (_T_839),	// matmul/matmul-hw.mlir:17821:13
    .p1_wr_en   (_T_843),	// matmul/matmul-hw.mlir:17808:13
    .p1_wr_data (_T_842),	// matmul/matmul-hw.mlir:17809:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2346)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3344 (	// matmul/matmul-hw.mlir:17655:36
    .p0_rd_en   (_T_834),	// matmul/matmul-hw.mlir:17851:13
    .p1_wr_en   (_T_838),	// matmul/matmul-hw.mlir:17838:13
    .p1_wr_data (_T_837),	// matmul/matmul-hw.mlir:17839:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2345)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3345 (	// matmul/matmul-hw.mlir:17656:36
    .p0_rd_en   (_T_829),	// matmul/matmul-hw.mlir:17881:13
    .p1_wr_en   (_T_833),	// matmul/matmul-hw.mlir:17868:13
    .p1_wr_data (_T_832),	// matmul/matmul-hw.mlir:17869:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2344)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3346 (	// matmul/matmul-hw.mlir:17657:36
    .p0_rd_en   (_T_824),	// matmul/matmul-hw.mlir:17911:13
    .p1_wr_en   (_T_828),	// matmul/matmul-hw.mlir:17898:13
    .p1_wr_data (_T_827),	// matmul/matmul-hw.mlir:17899:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2343)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3347 (	// matmul/matmul-hw.mlir:17658:36
    .p0_rd_en   (_T_819),	// matmul/matmul-hw.mlir:17941:13
    .p1_wr_en   (_T_823),	// matmul/matmul-hw.mlir:17928:13
    .p1_wr_data (_T_822),	// matmul/matmul-hw.mlir:17929:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2342)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3348 (	// matmul/matmul-hw.mlir:17659:37
    .p0_rd_en   (_T_814),	// matmul/matmul-hw.mlir:17971:13
    .p1_wr_en   (_T_818),	// matmul/matmul-hw.mlir:17958:13
    .p1_wr_data (_T_817),	// matmul/matmul-hw.mlir:17959:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2341)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3349 (	// matmul/matmul-hw.mlir:17660:37
    .p0_rd_en   (_T_809),	// matmul/matmul-hw.mlir:18001:13
    .p1_wr_en   (_T_813),	// matmul/matmul-hw.mlir:17988:13
    .p1_wr_data (_T_812),	// matmul/matmul-hw.mlir:17989:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2340)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3350 (	// matmul/matmul-hw.mlir:17661:37
    .p0_rd_en   (_T_804),	// matmul/matmul-hw.mlir:18031:13
    .p1_wr_en   (_T_808),	// matmul/matmul-hw.mlir:18018:13
    .p1_wr_data (_T_807),	// matmul/matmul-hw.mlir:18019:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2339)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3351 (	// matmul/matmul-hw.mlir:17662:37
    .p0_rd_en   (_T_799),	// matmul/matmul-hw.mlir:18061:13
    .p1_wr_en   (_T_803),	// matmul/matmul-hw.mlir:18048:13
    .p1_wr_data (_T_802),	// matmul/matmul-hw.mlir:18049:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2338)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3352 (	// matmul/matmul-hw.mlir:17663:37
    .p0_rd_en   (_T_794),	// matmul/matmul-hw.mlir:18091:13
    .p1_wr_en   (_T_798),	// matmul/matmul-hw.mlir:18078:13
    .p1_wr_data (_T_797),	// matmul/matmul-hw.mlir:18079:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2337)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3353 (	// matmul/matmul-hw.mlir:17664:37
    .p0_rd_en   (_T_789),	// matmul/matmul-hw.mlir:18121:13
    .p1_wr_en   (_T_793),	// matmul/matmul-hw.mlir:18108:13
    .p1_wr_data (_T_792),	// matmul/matmul-hw.mlir:18109:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2336)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3354 (	// matmul/matmul-hw.mlir:17665:37
    .p0_rd_en   (_T_786),	// matmul/matmul-hw.mlir:18148:13
    .p1_wr_en   (_T_788),	// matmul/matmul-hw.mlir:18138:13
    .p1_wr_data (_T_787),	// matmul/matmul-hw.mlir:18139:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2335)
  );
  assign _T_868 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17666:13
  assign _T_867 = _T_2808 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8902:19, :17667:13
  assign _T_866 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17668:13
  assign _T_865 = _T_2797 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17669:13
  mult mult_inst96 (	// matmul/matmul-hw.mlir:17670:27
    .a      (A_reg_bank96_p0_rd_data),	// matmul/matmul-hw.mlir:12311:32
    .b      (_T_2460),
    .t      (_T_2797),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst96_result)
  );
  assign _T_864 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17671:13
  assign a_i_k_0_i_j_6 = A_reg_bank96_p0_rd_data;	// matmul/matmul-hw.mlir:12311:32, :17673:5
  //PROBE: a_i_k_0_i_j_6	// matmul/matmul-hw.mlir:17674:5
  assign b_i_k_0_i_j_6 = _T_2460;	// matmul/matmul-hw.mlir:17676:5
  //PROBE: b_i_k_0_i_j_6	// matmul/matmul-hw.mlir:17677:5
  assign c_prev_i_k_0_i_j_6 = C_reg_bank0_p0_rd_data_2351;	// matmul/matmul-hw.mlir:17649:36, :17679:5
  //PROBE: c_prev_i_k_0_i_j_6	// matmul/matmul-hw.mlir:17680:5
  assign tk_i_k_0_i_j_6 = _T_2775;	// matmul/matmul-hw.mlir:17682:5
  //PROBE: tk_i_k_0_i_j_6	// matmul/matmul-hw.mlir:17683:5
  wire [31:0] _T_3355 = mult_inst96_result + C_reg_bank0_p0_rd_data_2351;	// matmul/matmul-hw.mlir:17649:36, :17670:27, :17684:13
  assign c_i_k_0_i_j_6 = _T_3355;	// matmul/matmul-hw.mlir:17686:5
  //PROBE: c_i_k_0_i_j_6	// matmul/matmul-hw.mlir:17687:5
  assign _T_863 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17688:13
  assign _T_862 = _T_2819 ? _T_3355 : 32'bx;	// matmul/matmul-hw.mlir:8897:19, :17689:13
  localparam [3:0] _T_3357 = 4'h0;	// matmul/matmul-hw.mlir:17692:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17693:5
    if (rst)	// matmul/matmul-hw.mlir:17693:5
      i_k_next_3356 <= _T_3357;	// matmul/matmul-hw.mlir:17696:7
    else	// matmul/matmul-hw.mlir:17693:5
      i_k_next_3356 <= i_j_next_3336;	// matmul/matmul-hw.mlir:17574:13, :17694:7
  end // always @(posedge)
  assign _T_861 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17698:13
  assign _T_860 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17699:13
  mult mult_inst97 (	// matmul/matmul-hw.mlir:17700:27
    .a      (A_reg_bank97_p0_rd_data),	// matmul/matmul-hw.mlir:12312:32
    .b      (_T_2476),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst97_result)
  );
  assign _T_859 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17701:13
  assign a_i_k_1_i_j_6 = A_reg_bank97_p0_rd_data;	// matmul/matmul-hw.mlir:12312:32, :17703:5
  //PROBE: a_i_k_1_i_j_6	// matmul/matmul-hw.mlir:17704:5
  assign b_i_k_1_i_j_6 = _T_2476;	// matmul/matmul-hw.mlir:17706:5
  //PROBE: b_i_k_1_i_j_6	// matmul/matmul-hw.mlir:17707:5
  assign c_prev_i_k_1_i_j_6 = C_reg_bank1_p0_rd_data_2350;	// matmul/matmul-hw.mlir:17650:36, :17709:5
  //PROBE: c_prev_i_k_1_i_j_6	// matmul/matmul-hw.mlir:17710:5
  assign tk_i_k_1_i_j_6 = _T_2786;	// matmul/matmul-hw.mlir:17712:5
  //PROBE: tk_i_k_1_i_j_6	// matmul/matmul-hw.mlir:17713:5
  wire [31:0] _T_3358 = mult_inst97_result + C_reg_bank1_p0_rd_data_2350;	// matmul/matmul-hw.mlir:17650:36, :17700:27, :17714:13
  assign c_i_k_1_i_j_6 = _T_3358;	// matmul/matmul-hw.mlir:17716:5
  //PROBE: c_i_k_1_i_j_6	// matmul/matmul-hw.mlir:17717:5
  assign _T_858 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17718:13
  assign _T_857 = _T_2830 ? _T_3358 : 32'bx;	// matmul/matmul-hw.mlir:8892:19, :17719:13
  localparam [3:0] _T_3360 = 4'h0;	// matmul/matmul-hw.mlir:17722:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17723:5
    if (rst)	// matmul/matmul-hw.mlir:17723:5
      i_k_next_3359 <= _T_3360;	// matmul/matmul-hw.mlir:17726:7
    else	// matmul/matmul-hw.mlir:17723:5
      i_k_next_3359 <= i_k_next_3356;	// matmul/matmul-hw.mlir:17691:13, :17724:7
  end // always @(posedge)
  assign _T_856 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17728:13
  assign _T_855 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17729:13
  mult mult_inst98 (	// matmul/matmul-hw.mlir:17730:27
    .a      (A_reg_bank98_p0_rd_data),	// matmul/matmul-hw.mlir:12313:32
    .b      (_T_2492),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst98_result)
  );
  assign _T_854 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17731:13
  assign a_i_k_2_i_j_6 = A_reg_bank98_p0_rd_data;	// matmul/matmul-hw.mlir:12313:32, :17733:5
  //PROBE: a_i_k_2_i_j_6	// matmul/matmul-hw.mlir:17734:5
  assign b_i_k_2_i_j_6 = _T_2492;	// matmul/matmul-hw.mlir:17736:5
  //PROBE: b_i_k_2_i_j_6	// matmul/matmul-hw.mlir:17737:5
  assign c_prev_i_k_2_i_j_6 = C_reg_bank2_p0_rd_data_2349;	// matmul/matmul-hw.mlir:17651:36, :17739:5
  //PROBE: c_prev_i_k_2_i_j_6	// matmul/matmul-hw.mlir:17740:5
  assign tk_i_k_2_i_j_6 = _T_2797;	// matmul/matmul-hw.mlir:17742:5
  //PROBE: tk_i_k_2_i_j_6	// matmul/matmul-hw.mlir:17743:5
  wire [31:0] _T_3361 = mult_inst98_result + C_reg_bank2_p0_rd_data_2349;	// matmul/matmul-hw.mlir:17651:36, :17730:27, :17744:13
  assign c_i_k_2_i_j_6 = _T_3361;	// matmul/matmul-hw.mlir:17746:5
  //PROBE: c_i_k_2_i_j_6	// matmul/matmul-hw.mlir:17747:5
  assign _T_853 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17748:13
  assign _T_852 = _T_2841 ? _T_3361 : 32'bx;	// matmul/matmul-hw.mlir:8887:19, :17749:13
  localparam [3:0] _T_3363 = 4'h0;	// matmul/matmul-hw.mlir:17752:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17753:5
    if (rst)	// matmul/matmul-hw.mlir:17753:5
      i_k_next_3362 <= _T_3363;	// matmul/matmul-hw.mlir:17756:7
    else	// matmul/matmul-hw.mlir:17753:5
      i_k_next_3362 <= i_k_next_3359;	// matmul/matmul-hw.mlir:17721:13, :17754:7
  end // always @(posedge)
  assign _T_851 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17758:13
  assign _T_850 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17759:13
  mult mult_inst99 (	// matmul/matmul-hw.mlir:17760:27
    .a      (A_reg_bank99_p0_rd_data),	// matmul/matmul-hw.mlir:12314:32
    .b      (_T_2508),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst99_result)
  );
  assign _T_849 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17761:13
  assign a_i_k_3_i_j_6 = A_reg_bank99_p0_rd_data;	// matmul/matmul-hw.mlir:12314:32, :17763:5
  //PROBE: a_i_k_3_i_j_6	// matmul/matmul-hw.mlir:17764:5
  assign b_i_k_3_i_j_6 = _T_2508;	// matmul/matmul-hw.mlir:17766:5
  //PROBE: b_i_k_3_i_j_6	// matmul/matmul-hw.mlir:17767:5
  assign c_prev_i_k_3_i_j_6 = C_reg_bank3_p0_rd_data_2348;	// matmul/matmul-hw.mlir:17652:36, :17769:5
  //PROBE: c_prev_i_k_3_i_j_6	// matmul/matmul-hw.mlir:17770:5
  assign tk_i_k_3_i_j_6 = _T_2808;	// matmul/matmul-hw.mlir:17772:5
  //PROBE: tk_i_k_3_i_j_6	// matmul/matmul-hw.mlir:17773:5
  wire [31:0] _T_3364 = mult_inst99_result + C_reg_bank3_p0_rd_data_2348;	// matmul/matmul-hw.mlir:17652:36, :17760:27, :17774:13
  assign c_i_k_3_i_j_6 = _T_3364;	// matmul/matmul-hw.mlir:17776:5
  //PROBE: c_i_k_3_i_j_6	// matmul/matmul-hw.mlir:17777:5
  assign _T_848 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17778:13
  assign _T_847 = _T_2852 ? _T_3364 : 32'bx;	// matmul/matmul-hw.mlir:8882:19, :17779:13
  localparam [3:0] _T_3366 = 4'h0;	// matmul/matmul-hw.mlir:17782:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17783:5
    if (rst)	// matmul/matmul-hw.mlir:17783:5
      i_k_next_3365 <= _T_3366;	// matmul/matmul-hw.mlir:17786:7
    else	// matmul/matmul-hw.mlir:17783:5
      i_k_next_3365 <= i_k_next_3362;	// matmul/matmul-hw.mlir:17751:13, :17784:7
  end // always @(posedge)
  assign _T_846 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17788:13
  assign _T_845 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17789:13
  mult mult_inst100 (	// matmul/matmul-hw.mlir:17790:28
    .a      (A_reg_bank100_p0_rd_data),	// matmul/matmul-hw.mlir:12315:33
    .b      (_T_2524),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst100_result)
  );
  assign _T_844 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17791:13
  assign a_i_k_4_i_j_6 = A_reg_bank100_p0_rd_data;	// matmul/matmul-hw.mlir:12315:33, :17793:5
  //PROBE: a_i_k_4_i_j_6	// matmul/matmul-hw.mlir:17794:5
  assign b_i_k_4_i_j_6 = _T_2524;	// matmul/matmul-hw.mlir:17796:5
  //PROBE: b_i_k_4_i_j_6	// matmul/matmul-hw.mlir:17797:5
  assign c_prev_i_k_4_i_j_6 = C_reg_bank4_p0_rd_data_2347;	// matmul/matmul-hw.mlir:17653:36, :17799:5
  //PROBE: c_prev_i_k_4_i_j_6	// matmul/matmul-hw.mlir:17800:5
  assign tk_i_k_4_i_j_6 = _T_2819;	// matmul/matmul-hw.mlir:17802:5
  //PROBE: tk_i_k_4_i_j_6	// matmul/matmul-hw.mlir:17803:5
  wire [31:0] _T_3367 = mult_inst100_result + C_reg_bank4_p0_rd_data_2347;	// matmul/matmul-hw.mlir:17653:36, :17790:28, :17804:13
  assign c_i_k_4_i_j_6 = _T_3367;	// matmul/matmul-hw.mlir:17806:5
  //PROBE: c_i_k_4_i_j_6	// matmul/matmul-hw.mlir:17807:5
  assign _T_843 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17808:13
  assign _T_842 = _T_2863 ? _T_3367 : 32'bx;	// matmul/matmul-hw.mlir:8877:19, :17809:13
  localparam [3:0] _T_3369 = 4'h0;	// matmul/matmul-hw.mlir:17812:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17813:5
    if (rst)	// matmul/matmul-hw.mlir:17813:5
      i_k_next_3368 <= _T_3369;	// matmul/matmul-hw.mlir:17816:7
    else	// matmul/matmul-hw.mlir:17813:5
      i_k_next_3368 <= i_k_next_3365;	// matmul/matmul-hw.mlir:17781:13, :17814:7
  end // always @(posedge)
  assign _T_841 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17818:13
  assign _T_840 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17819:13
  mult mult_inst101 (	// matmul/matmul-hw.mlir:17820:28
    .a      (A_reg_bank101_p0_rd_data),	// matmul/matmul-hw.mlir:12316:33
    .b      (_T_2540),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst101_result)
  );
  assign _T_839 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17821:13
  assign a_i_k_5_i_j_6 = A_reg_bank101_p0_rd_data;	// matmul/matmul-hw.mlir:12316:33, :17823:5
  //PROBE: a_i_k_5_i_j_6	// matmul/matmul-hw.mlir:17824:5
  assign b_i_k_5_i_j_6 = _T_2540;	// matmul/matmul-hw.mlir:17826:5
  //PROBE: b_i_k_5_i_j_6	// matmul/matmul-hw.mlir:17827:5
  assign c_prev_i_k_5_i_j_6 = C_reg_bank5_p0_rd_data_2346;	// matmul/matmul-hw.mlir:17654:36, :17829:5
  //PROBE: c_prev_i_k_5_i_j_6	// matmul/matmul-hw.mlir:17830:5
  assign tk_i_k_5_i_j_6 = _T_2830;	// matmul/matmul-hw.mlir:17832:5
  //PROBE: tk_i_k_5_i_j_6	// matmul/matmul-hw.mlir:17833:5
  wire [31:0] _T_3370 = mult_inst101_result + C_reg_bank5_p0_rd_data_2346;	// matmul/matmul-hw.mlir:17654:36, :17820:28, :17834:13
  assign c_i_k_5_i_j_6 = _T_3370;	// matmul/matmul-hw.mlir:17836:5
  //PROBE: c_i_k_5_i_j_6	// matmul/matmul-hw.mlir:17837:5
  assign _T_838 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17838:13
  assign _T_837 = _T_2874 ? _T_3370 : 32'bx;	// matmul/matmul-hw.mlir:8872:19, :17839:13
  localparam [3:0] _T_3372 = 4'h0;	// matmul/matmul-hw.mlir:17842:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17843:5
    if (rst)	// matmul/matmul-hw.mlir:17843:5
      i_k_next_3371 <= _T_3372;	// matmul/matmul-hw.mlir:17846:7
    else	// matmul/matmul-hw.mlir:17843:5
      i_k_next_3371 <= i_k_next_3368;	// matmul/matmul-hw.mlir:17811:13, :17844:7
  end // always @(posedge)
  assign _T_836 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17848:13
  assign _T_835 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17849:13
  mult mult_inst102 (	// matmul/matmul-hw.mlir:17850:28
    .a      (A_reg_bank102_p0_rd_data),	// matmul/matmul-hw.mlir:12317:33
    .b      (_T_2556),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst102_result)
  );
  assign _T_834 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17851:13
  assign a_i_k_6_i_j_6 = A_reg_bank102_p0_rd_data;	// matmul/matmul-hw.mlir:12317:33, :17853:5
  //PROBE: a_i_k_6_i_j_6	// matmul/matmul-hw.mlir:17854:5
  assign b_i_k_6_i_j_6 = _T_2556;	// matmul/matmul-hw.mlir:17856:5
  //PROBE: b_i_k_6_i_j_6	// matmul/matmul-hw.mlir:17857:5
  assign c_prev_i_k_6_i_j_6 = C_reg_bank6_p0_rd_data_2345;	// matmul/matmul-hw.mlir:17655:36, :17859:5
  //PROBE: c_prev_i_k_6_i_j_6	// matmul/matmul-hw.mlir:17860:5
  assign tk_i_k_6_i_j_6 = _T_2841;	// matmul/matmul-hw.mlir:17862:5
  //PROBE: tk_i_k_6_i_j_6	// matmul/matmul-hw.mlir:17863:5
  wire [31:0] _T_3373 = mult_inst102_result + C_reg_bank6_p0_rd_data_2345;	// matmul/matmul-hw.mlir:17655:36, :17850:28, :17864:13
  assign c_i_k_6_i_j_6 = _T_3373;	// matmul/matmul-hw.mlir:17866:5
  //PROBE: c_i_k_6_i_j_6	// matmul/matmul-hw.mlir:17867:5
  assign _T_833 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17868:13
  assign _T_832 = _T_2885 ? _T_3373 : 32'bx;	// matmul/matmul-hw.mlir:8867:19, :17869:13
  localparam [3:0] _T_3375 = 4'h0;	// matmul/matmul-hw.mlir:17872:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17873:5
    if (rst)	// matmul/matmul-hw.mlir:17873:5
      i_k_next_3374 <= _T_3375;	// matmul/matmul-hw.mlir:17876:7
    else	// matmul/matmul-hw.mlir:17873:5
      i_k_next_3374 <= i_k_next_3371;	// matmul/matmul-hw.mlir:17841:13, :17874:7
  end // always @(posedge)
  assign _T_831 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17878:13
  assign _T_830 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17879:13
  mult mult_inst103 (	// matmul/matmul-hw.mlir:17880:28
    .a      (A_reg_bank103_p0_rd_data),	// matmul/matmul-hw.mlir:12318:33
    .b      (_T_2572),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst103_result)
  );
  assign _T_829 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17881:13
  assign a_i_k_7_i_j_6 = A_reg_bank103_p0_rd_data;	// matmul/matmul-hw.mlir:12318:33, :17883:5
  //PROBE: a_i_k_7_i_j_6	// matmul/matmul-hw.mlir:17884:5
  assign b_i_k_7_i_j_6 = _T_2572;	// matmul/matmul-hw.mlir:17886:5
  //PROBE: b_i_k_7_i_j_6	// matmul/matmul-hw.mlir:17887:5
  assign c_prev_i_k_7_i_j_6 = C_reg_bank7_p0_rd_data_2344;	// matmul/matmul-hw.mlir:17656:36, :17889:5
  //PROBE: c_prev_i_k_7_i_j_6	// matmul/matmul-hw.mlir:17890:5
  assign tk_i_k_7_i_j_6 = _T_2852;	// matmul/matmul-hw.mlir:17892:5
  //PROBE: tk_i_k_7_i_j_6	// matmul/matmul-hw.mlir:17893:5
  wire [31:0] _T_3376 = mult_inst103_result + C_reg_bank7_p0_rd_data_2344;	// matmul/matmul-hw.mlir:17656:36, :17880:28, :17894:13
  assign c_i_k_7_i_j_6 = _T_3376;	// matmul/matmul-hw.mlir:17896:5
  //PROBE: c_i_k_7_i_j_6	// matmul/matmul-hw.mlir:17897:5
  assign _T_828 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17898:13
  assign _T_827 = _T_2892 ? _T_3376 : 32'bx;	// matmul/matmul-hw.mlir:8862:19, :17899:13
  localparam [3:0] _T_3378 = 4'h0;	// matmul/matmul-hw.mlir:17902:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17903:5
    if (rst)	// matmul/matmul-hw.mlir:17903:5
      i_k_next_3377 <= _T_3378;	// matmul/matmul-hw.mlir:17906:7
    else	// matmul/matmul-hw.mlir:17903:5
      i_k_next_3377 <= i_k_next_3374;	// matmul/matmul-hw.mlir:17871:13, :17904:7
  end // always @(posedge)
  assign _T_826 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17908:13
  assign _T_825 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17909:13
  mult mult_inst104 (	// matmul/matmul-hw.mlir:17910:28
    .a      (A_reg_bank104_p0_rd_data),	// matmul/matmul-hw.mlir:12319:33
    .b      (_T_2588),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst104_result)
  );
  assign _T_824 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17911:13
  assign a_i_k_8_i_j_6 = A_reg_bank104_p0_rd_data;	// matmul/matmul-hw.mlir:12319:33, :17913:5
  //PROBE: a_i_k_8_i_j_6	// matmul/matmul-hw.mlir:17914:5
  assign b_i_k_8_i_j_6 = _T_2588;	// matmul/matmul-hw.mlir:17916:5
  //PROBE: b_i_k_8_i_j_6	// matmul/matmul-hw.mlir:17917:5
  assign c_prev_i_k_8_i_j_6 = C_reg_bank8_p0_rd_data_2343;	// matmul/matmul-hw.mlir:17657:36, :17919:5
  //PROBE: c_prev_i_k_8_i_j_6	// matmul/matmul-hw.mlir:17920:5
  assign tk_i_k_8_i_j_6 = _T_2863;	// matmul/matmul-hw.mlir:17922:5
  //PROBE: tk_i_k_8_i_j_6	// matmul/matmul-hw.mlir:17923:5
  wire [31:0] _T_3379 = mult_inst104_result + C_reg_bank8_p0_rd_data_2343;	// matmul/matmul-hw.mlir:17657:36, :17910:28, :17924:13
  assign c_i_k_8_i_j_6 = _T_3379;	// matmul/matmul-hw.mlir:17926:5
  //PROBE: c_i_k_8_i_j_6	// matmul/matmul-hw.mlir:17927:5
  assign _T_823 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17928:13
  assign _T_822 = _T_2897 ? _T_3379 : 32'bx;	// matmul/matmul-hw.mlir:8857:19, :17929:13
  localparam [3:0] _T_3381 = 4'h0;	// matmul/matmul-hw.mlir:17932:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17933:5
    if (rst)	// matmul/matmul-hw.mlir:17933:5
      i_k_next_3380 <= _T_3381;	// matmul/matmul-hw.mlir:17936:7
    else	// matmul/matmul-hw.mlir:17933:5
      i_k_next_3380 <= i_k_next_3377;	// matmul/matmul-hw.mlir:17901:13, :17934:7
  end // always @(posedge)
  assign _T_821 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17938:13
  assign _T_820 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17939:13
  mult mult_inst105 (	// matmul/matmul-hw.mlir:17940:28
    .a      (A_reg_bank105_p0_rd_data),	// matmul/matmul-hw.mlir:12320:33
    .b      (_T_2604),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst105_result)
  );
  assign _T_819 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17941:13
  assign a_i_k_9_i_j_6 = A_reg_bank105_p0_rd_data;	// matmul/matmul-hw.mlir:12320:33, :17943:5
  //PROBE: a_i_k_9_i_j_6	// matmul/matmul-hw.mlir:17944:5
  assign b_i_k_9_i_j_6 = _T_2604;	// matmul/matmul-hw.mlir:17946:5
  //PROBE: b_i_k_9_i_j_6	// matmul/matmul-hw.mlir:17947:5
  assign c_prev_i_k_9_i_j_6 = C_reg_bank9_p0_rd_data_2342;	// matmul/matmul-hw.mlir:17658:36, :17949:5
  //PROBE: c_prev_i_k_9_i_j_6	// matmul/matmul-hw.mlir:17950:5
  assign tk_i_k_9_i_j_6 = _T_2874;	// matmul/matmul-hw.mlir:17952:5
  //PROBE: tk_i_k_9_i_j_6	// matmul/matmul-hw.mlir:17953:5
  wire [31:0] _T_3382 = mult_inst105_result + C_reg_bank9_p0_rd_data_2342;	// matmul/matmul-hw.mlir:17658:36, :17940:28, :17954:13
  assign c_i_k_9_i_j_6 = _T_3382;	// matmul/matmul-hw.mlir:17956:5
  //PROBE: c_i_k_9_i_j_6	// matmul/matmul-hw.mlir:17957:5
  assign _T_818 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17958:13
  assign _T_817 = _T_2902 ? _T_3382 : 32'bx;	// matmul/matmul-hw.mlir:8852:19, :17959:13
  localparam [3:0] _T_3384 = 4'h0;	// matmul/matmul-hw.mlir:17962:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17963:5
    if (rst)	// matmul/matmul-hw.mlir:17963:5
      i_k_next_3383 <= _T_3384;	// matmul/matmul-hw.mlir:17966:7
    else	// matmul/matmul-hw.mlir:17963:5
      i_k_next_3383 <= i_k_next_3380;	// matmul/matmul-hw.mlir:17931:13, :17964:7
  end // always @(posedge)
  assign _T_816 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17968:13
  assign _T_815 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17969:13
  mult mult_inst106 (	// matmul/matmul-hw.mlir:17970:28
    .a      (A_reg_bank106_p0_rd_data),	// matmul/matmul-hw.mlir:12321:33
    .b      (_T_2620),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst106_result)
  );
  assign _T_814 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17971:13
  assign a_i_k_10_i_j_6 = A_reg_bank106_p0_rd_data;	// matmul/matmul-hw.mlir:12321:33, :17973:5
  //PROBE: a_i_k_10_i_j_6	// matmul/matmul-hw.mlir:17974:5
  assign b_i_k_10_i_j_6 = _T_2620;	// matmul/matmul-hw.mlir:17976:5
  //PROBE: b_i_k_10_i_j_6	// matmul/matmul-hw.mlir:17977:5
  assign c_prev_i_k_10_i_j_6 = C_reg_bank10_p0_rd_data_2341;	// matmul/matmul-hw.mlir:17659:37, :17979:5
  //PROBE: c_prev_i_k_10_i_j_6	// matmul/matmul-hw.mlir:17980:5
  assign tk_i_k_10_i_j_6 = _T_2885;	// matmul/matmul-hw.mlir:17982:5
  //PROBE: tk_i_k_10_i_j_6	// matmul/matmul-hw.mlir:17983:5
  wire [31:0] _T_3385 = mult_inst106_result + C_reg_bank10_p0_rd_data_2341;	// matmul/matmul-hw.mlir:17659:37, :17970:28, :17984:13
  assign c_i_k_10_i_j_6 = _T_3385;	// matmul/matmul-hw.mlir:17986:5
  //PROBE: c_i_k_10_i_j_6	// matmul/matmul-hw.mlir:17987:5
  assign _T_813 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17988:13
  assign _T_812 = _T_2907 ? _T_3385 : 32'bx;	// matmul/matmul-hw.mlir:8847:19, :17989:13
  localparam [3:0] _T_3387 = 4'h0;	// matmul/matmul-hw.mlir:17992:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:17993:5
    if (rst)	// matmul/matmul-hw.mlir:17993:5
      i_k_next_3386 <= _T_3387;	// matmul/matmul-hw.mlir:17996:7
    else	// matmul/matmul-hw.mlir:17993:5
      i_k_next_3386 <= i_k_next_3383;	// matmul/matmul-hw.mlir:17961:13, :17994:7
  end // always @(posedge)
  assign _T_811 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17998:13
  assign _T_810 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :17999:13
  mult mult_inst107 (	// matmul/matmul-hw.mlir:18000:28
    .a      (A_reg_bank107_p0_rd_data),	// matmul/matmul-hw.mlir:12322:33
    .b      (_T_2636),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst107_result)
  );
  assign _T_809 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18001:13
  assign a_i_k_11_i_j_6 = A_reg_bank107_p0_rd_data;	// matmul/matmul-hw.mlir:12322:33, :18003:5
  //PROBE: a_i_k_11_i_j_6	// matmul/matmul-hw.mlir:18004:5
  assign b_i_k_11_i_j_6 = _T_2636;	// matmul/matmul-hw.mlir:18006:5
  //PROBE: b_i_k_11_i_j_6	// matmul/matmul-hw.mlir:18007:5
  assign c_prev_i_k_11_i_j_6 = C_reg_bank11_p0_rd_data_2340;	// matmul/matmul-hw.mlir:17660:37, :18009:5
  //PROBE: c_prev_i_k_11_i_j_6	// matmul/matmul-hw.mlir:18010:5
  assign tk_i_k_11_i_j_6 = _T_2892;	// matmul/matmul-hw.mlir:18012:5
  //PROBE: tk_i_k_11_i_j_6	// matmul/matmul-hw.mlir:18013:5
  wire [31:0] _T_3388 = mult_inst107_result + C_reg_bank11_p0_rd_data_2340;	// matmul/matmul-hw.mlir:17660:37, :18000:28, :18014:13
  assign c_i_k_11_i_j_6 = _T_3388;	// matmul/matmul-hw.mlir:18016:5
  //PROBE: c_i_k_11_i_j_6	// matmul/matmul-hw.mlir:18017:5
  assign _T_808 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18018:13
  assign _T_807 = _T_2912 ? _T_3388 : 32'bx;	// matmul/matmul-hw.mlir:8842:19, :18019:13
  localparam [3:0] _T_3390 = 4'h0;	// matmul/matmul-hw.mlir:18022:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18023:5
    if (rst)	// matmul/matmul-hw.mlir:18023:5
      i_k_next_3389 <= _T_3390;	// matmul/matmul-hw.mlir:18026:7
    else	// matmul/matmul-hw.mlir:18023:5
      i_k_next_3389 <= i_k_next_3386;	// matmul/matmul-hw.mlir:17991:13, :18024:7
  end // always @(posedge)
  assign _T_806 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18028:13
  assign _T_805 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18029:13
  mult mult_inst108 (	// matmul/matmul-hw.mlir:18030:28
    .a      (A_reg_bank108_p0_rd_data),	// matmul/matmul-hw.mlir:12323:33
    .b      (_T_2652),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst108_result)
  );
  assign _T_804 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18031:13
  assign a_i_k_12_i_j_6 = A_reg_bank108_p0_rd_data;	// matmul/matmul-hw.mlir:12323:33, :18033:5
  //PROBE: a_i_k_12_i_j_6	// matmul/matmul-hw.mlir:18034:5
  assign b_i_k_12_i_j_6 = _T_2652;	// matmul/matmul-hw.mlir:18036:5
  //PROBE: b_i_k_12_i_j_6	// matmul/matmul-hw.mlir:18037:5
  assign c_prev_i_k_12_i_j_6 = C_reg_bank12_p0_rd_data_2339;	// matmul/matmul-hw.mlir:17661:37, :18039:5
  //PROBE: c_prev_i_k_12_i_j_6	// matmul/matmul-hw.mlir:18040:5
  assign tk_i_k_12_i_j_6 = _T_2897;	// matmul/matmul-hw.mlir:18042:5
  //PROBE: tk_i_k_12_i_j_6	// matmul/matmul-hw.mlir:18043:5
  wire [31:0] _T_3391 = mult_inst108_result + C_reg_bank12_p0_rd_data_2339;	// matmul/matmul-hw.mlir:17661:37, :18030:28, :18044:13
  assign c_i_k_12_i_j_6 = _T_3391;	// matmul/matmul-hw.mlir:18046:5
  //PROBE: c_i_k_12_i_j_6	// matmul/matmul-hw.mlir:18047:5
  assign _T_803 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18048:13
  assign _T_802 = _T_2917 ? _T_3391 : 32'bx;	// matmul/matmul-hw.mlir:8837:19, :18049:13
  localparam [3:0] _T_3393 = 4'h0;	// matmul/matmul-hw.mlir:18052:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18053:5
    if (rst)	// matmul/matmul-hw.mlir:18053:5
      i_k_next_3392 <= _T_3393;	// matmul/matmul-hw.mlir:18056:7
    else	// matmul/matmul-hw.mlir:18053:5
      i_k_next_3392 <= i_k_next_3389;	// matmul/matmul-hw.mlir:18021:13, :18054:7
  end // always @(posedge)
  assign _T_801 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18058:13
  assign _T_800 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18059:13
  mult mult_inst109 (	// matmul/matmul-hw.mlir:18060:28
    .a      (A_reg_bank109_p0_rd_data),	// matmul/matmul-hw.mlir:12324:33
    .b      (_T_2668),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst109_result)
  );
  assign _T_799 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18061:13
  assign a_i_k_13_i_j_6 = A_reg_bank109_p0_rd_data;	// matmul/matmul-hw.mlir:12324:33, :18063:5
  //PROBE: a_i_k_13_i_j_6	// matmul/matmul-hw.mlir:18064:5
  assign b_i_k_13_i_j_6 = _T_2668;	// matmul/matmul-hw.mlir:18066:5
  //PROBE: b_i_k_13_i_j_6	// matmul/matmul-hw.mlir:18067:5
  assign c_prev_i_k_13_i_j_6 = C_reg_bank13_p0_rd_data_2338;	// matmul/matmul-hw.mlir:17662:37, :18069:5
  //PROBE: c_prev_i_k_13_i_j_6	// matmul/matmul-hw.mlir:18070:5
  assign tk_i_k_13_i_j_6 = _T_2902;	// matmul/matmul-hw.mlir:18072:5
  //PROBE: tk_i_k_13_i_j_6	// matmul/matmul-hw.mlir:18073:5
  wire [31:0] _T_3394 = mult_inst109_result + C_reg_bank13_p0_rd_data_2338;	// matmul/matmul-hw.mlir:17662:37, :18060:28, :18074:13
  assign c_i_k_13_i_j_6 = _T_3394;	// matmul/matmul-hw.mlir:18076:5
  //PROBE: c_i_k_13_i_j_6	// matmul/matmul-hw.mlir:18077:5
  assign _T_798 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18078:13
  assign _T_797 = _T_2922 ? _T_3394 : 32'bx;	// matmul/matmul-hw.mlir:8832:19, :18079:13
  localparam [3:0] _T_3396 = 4'h0;	// matmul/matmul-hw.mlir:18082:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18083:5
    if (rst)	// matmul/matmul-hw.mlir:18083:5
      i_k_next_3395 <= _T_3396;	// matmul/matmul-hw.mlir:18086:7
    else	// matmul/matmul-hw.mlir:18083:5
      i_k_next_3395 <= i_k_next_3392;	// matmul/matmul-hw.mlir:18051:13, :18084:7
  end // always @(posedge)
  assign _T_796 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18088:13
  assign _T_795 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18089:13
  mult mult_inst110 (	// matmul/matmul-hw.mlir:18090:28
    .a      (A_reg_bank110_p0_rd_data),	// matmul/matmul-hw.mlir:12325:33
    .b      (_T_2684),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst110_result)
  );
  assign _T_794 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18091:13
  assign a_i_k_14_i_j_6 = A_reg_bank110_p0_rd_data;	// matmul/matmul-hw.mlir:12325:33, :18093:5
  //PROBE: a_i_k_14_i_j_6	// matmul/matmul-hw.mlir:18094:5
  assign b_i_k_14_i_j_6 = _T_2684;	// matmul/matmul-hw.mlir:18096:5
  //PROBE: b_i_k_14_i_j_6	// matmul/matmul-hw.mlir:18097:5
  assign c_prev_i_k_14_i_j_6 = C_reg_bank14_p0_rd_data_2337;	// matmul/matmul-hw.mlir:17663:37, :18099:5
  //PROBE: c_prev_i_k_14_i_j_6	// matmul/matmul-hw.mlir:18100:5
  assign tk_i_k_14_i_j_6 = _T_2907;	// matmul/matmul-hw.mlir:18102:5
  //PROBE: tk_i_k_14_i_j_6	// matmul/matmul-hw.mlir:18103:5
  wire [31:0] _T_3397 = mult_inst110_result + C_reg_bank14_p0_rd_data_2337;	// matmul/matmul-hw.mlir:17663:37, :18090:28, :18104:13
  assign c_i_k_14_i_j_6 = _T_3397;	// matmul/matmul-hw.mlir:18106:5
  //PROBE: c_i_k_14_i_j_6	// matmul/matmul-hw.mlir:18107:5
  assign _T_793 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18108:13
  assign _T_792 = _T_2927 ? _T_3397 : 32'bx;	// matmul/matmul-hw.mlir:8827:19, :18109:13
  localparam [3:0] _T_3399 = 4'h0;	// matmul/matmul-hw.mlir:18112:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18113:5
    if (rst)	// matmul/matmul-hw.mlir:18113:5
      i_k_next_3398 <= _T_3399;	// matmul/matmul-hw.mlir:18116:7
    else	// matmul/matmul-hw.mlir:18113:5
      i_k_next_3398 <= i_k_next_3395;	// matmul/matmul-hw.mlir:18081:13, :18114:7
  end // always @(posedge)
  assign _T_791 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18118:13
  assign _T_790 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18119:13
  mult mult_inst111 (	// matmul/matmul-hw.mlir:18120:28
    .a      (A_reg_bank111_p0_rd_data),	// matmul/matmul-hw.mlir:12326:33
    .b      (_T_2700),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst111_result)
  );
  assign _T_789 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18121:13
  assign a_i_k_15_i_j_6 = A_reg_bank111_p0_rd_data;	// matmul/matmul-hw.mlir:12326:33, :18123:5
  //PROBE: a_i_k_15_i_j_6	// matmul/matmul-hw.mlir:18124:5
  assign b_i_k_15_i_j_6 = _T_2700;	// matmul/matmul-hw.mlir:18126:5
  //PROBE: b_i_k_15_i_j_6	// matmul/matmul-hw.mlir:18127:5
  assign c_prev_i_k_15_i_j_6 = C_reg_bank15_p0_rd_data_2336;	// matmul/matmul-hw.mlir:17664:37, :18129:5
  //PROBE: c_prev_i_k_15_i_j_6	// matmul/matmul-hw.mlir:18130:5
  assign tk_i_k_15_i_j_6 = _T_2912;	// matmul/matmul-hw.mlir:18132:5
  //PROBE: tk_i_k_15_i_j_6	// matmul/matmul-hw.mlir:18133:5
  wire [31:0] _T_3400 = mult_inst111_result + C_reg_bank15_p0_rd_data_2336;	// matmul/matmul-hw.mlir:17664:37, :18120:28, :18134:13
  assign c_i_k_15_i_j_6 = _T_3400;	// matmul/matmul-hw.mlir:18136:5
  //PROBE: c_i_k_15_i_j_6	// matmul/matmul-hw.mlir:18137:5
  assign _T_788 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18138:13
  assign _T_787 = _T_2932 ? _T_3400 : 32'bx;	// matmul/matmul-hw.mlir:8822:19, :18139:13
  localparam [3:0] _T_3402 = 4'h0;	// matmul/matmul-hw.mlir:18142:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18143:5
    if (rst)	// matmul/matmul-hw.mlir:18143:5
      i_k_next_3401 <= _T_3402;	// matmul/matmul-hw.mlir:18146:7
    else	// matmul/matmul-hw.mlir:18143:5
      i_k_next_3401 <= i_k_next_3398;	// matmul/matmul-hw.mlir:18111:13, :18144:7
  end // always @(posedge)
  assign _T_786 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18148:13
  wire [3:0][3:0] _T_3404 = i_delayed_3403;	// matmul/matmul-hw.mlir:18150:13
  wire [3:0][3:0] _T_3405 = {_T_3404[2'h0+:3], {{i_k_next_3401}}};	// matmul/matmul-hw.mlir:18141:13, :18151:19, :18152:13, :18153:13, :18154:13
  wire [3:0][3:0] _T_3406 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:18155:19, :18156:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18157:5
    if (rst)	// matmul/matmul-hw.mlir:18157:5
      i_delayed_3403 <= _T_3406;	// matmul/matmul-hw.mlir:18160:7
    else	// matmul/matmul-hw.mlir:18157:5
      i_delayed_3403 <= _T_3405;	// matmul/matmul-hw.mlir:18158:7
  end // always @(posedge)
  assign _T_785 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18164:13
  assign _T_784 = _T_2937 ? i_delayed_3403[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8819:18, :18150:13, :18162:20, :18163:13, :18165:13
  assign _T_783 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18166:13
  assign _T_782 = _T_2937 ? C_reg_bank16_p0_rd_data_2335 : 32'bx;	// matmul/matmul-hw.mlir:8817:19, :17665:37, :18167:13
  localparam [3:0] _T_3408 = 4'h0;	// matmul/matmul-hw.mlir:18170:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18171:5
    if (rst)	// matmul/matmul-hw.mlir:18171:5
      i_j_next_3407 <= _T_3408;	// matmul/matmul-hw.mlir:18174:7
    else	// matmul/matmul-hw.mlir:18171:5
      i_j_next_3407 <= i_j_next_3336;	// matmul/matmul-hw.mlir:17574:13, :18172:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3409 (	// matmul/matmul-hw.mlir:18244:36
    .p0_rd_en   (_T_777),	// matmul/matmul-hw.mlir:18266:13
    .p1_wr_en   (_T_781),	// matmul/matmul-hw.mlir:18261:13
    .p1_wr_data (_T_780),	// matmul/matmul-hw.mlir:18262:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2334)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3410 (	// matmul/matmul-hw.mlir:18245:36
    .p0_rd_en   (_T_772),	// matmul/matmul-hw.mlir:18296:13
    .p1_wr_en   (_T_776),	// matmul/matmul-hw.mlir:18283:13
    .p1_wr_data (_T_775),	// matmul/matmul-hw.mlir:18284:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2333)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3411 (	// matmul/matmul-hw.mlir:18246:36
    .p0_rd_en   (_T_767),	// matmul/matmul-hw.mlir:18326:13
    .p1_wr_en   (_T_771),	// matmul/matmul-hw.mlir:18313:13
    .p1_wr_data (_T_770),	// matmul/matmul-hw.mlir:18314:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2332)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3412 (	// matmul/matmul-hw.mlir:18247:36
    .p0_rd_en   (_T_762),	// matmul/matmul-hw.mlir:18356:13
    .p1_wr_en   (_T_766),	// matmul/matmul-hw.mlir:18343:13
    .p1_wr_data (_T_765),	// matmul/matmul-hw.mlir:18344:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2331)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3413 (	// matmul/matmul-hw.mlir:18248:36
    .p0_rd_en   (_T_757),	// matmul/matmul-hw.mlir:18386:13
    .p1_wr_en   (_T_761),	// matmul/matmul-hw.mlir:18373:13
    .p1_wr_data (_T_760),	// matmul/matmul-hw.mlir:18374:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2330)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3414 (	// matmul/matmul-hw.mlir:18249:36
    .p0_rd_en   (_T_752),	// matmul/matmul-hw.mlir:18416:13
    .p1_wr_en   (_T_756),	// matmul/matmul-hw.mlir:18403:13
    .p1_wr_data (_T_755),	// matmul/matmul-hw.mlir:18404:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2329)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3415 (	// matmul/matmul-hw.mlir:18250:36
    .p0_rd_en   (_T_747),	// matmul/matmul-hw.mlir:18446:13
    .p1_wr_en   (_T_751),	// matmul/matmul-hw.mlir:18433:13
    .p1_wr_data (_T_750),	// matmul/matmul-hw.mlir:18434:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2328)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3416 (	// matmul/matmul-hw.mlir:18251:36
    .p0_rd_en   (_T_742),	// matmul/matmul-hw.mlir:18476:13
    .p1_wr_en   (_T_746),	// matmul/matmul-hw.mlir:18463:13
    .p1_wr_data (_T_745),	// matmul/matmul-hw.mlir:18464:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2327)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3417 (	// matmul/matmul-hw.mlir:18252:36
    .p0_rd_en   (_T_737),	// matmul/matmul-hw.mlir:18506:13
    .p1_wr_en   (_T_741),	// matmul/matmul-hw.mlir:18493:13
    .p1_wr_data (_T_740),	// matmul/matmul-hw.mlir:18494:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2326)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3418 (	// matmul/matmul-hw.mlir:18253:36
    .p0_rd_en   (_T_732),	// matmul/matmul-hw.mlir:18536:13
    .p1_wr_en   (_T_736),	// matmul/matmul-hw.mlir:18523:13
    .p1_wr_data (_T_735),	// matmul/matmul-hw.mlir:18524:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2325)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3419 (	// matmul/matmul-hw.mlir:18254:37
    .p0_rd_en   (_T_727),	// matmul/matmul-hw.mlir:18566:13
    .p1_wr_en   (_T_731),	// matmul/matmul-hw.mlir:18553:13
    .p1_wr_data (_T_730),	// matmul/matmul-hw.mlir:18554:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2324)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3420 (	// matmul/matmul-hw.mlir:18255:37
    .p0_rd_en   (_T_722),	// matmul/matmul-hw.mlir:18596:13
    .p1_wr_en   (_T_726),	// matmul/matmul-hw.mlir:18583:13
    .p1_wr_data (_T_725),	// matmul/matmul-hw.mlir:18584:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2323)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3421 (	// matmul/matmul-hw.mlir:18256:37
    .p0_rd_en   (_T_717),	// matmul/matmul-hw.mlir:18626:13
    .p1_wr_en   (_T_721),	// matmul/matmul-hw.mlir:18613:13
    .p1_wr_data (_T_720),	// matmul/matmul-hw.mlir:18614:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2322)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3422 (	// matmul/matmul-hw.mlir:18257:37
    .p0_rd_en   (_T_712),	// matmul/matmul-hw.mlir:18656:13
    .p1_wr_en   (_T_716),	// matmul/matmul-hw.mlir:18643:13
    .p1_wr_data (_T_715),	// matmul/matmul-hw.mlir:18644:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2321)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3423 (	// matmul/matmul-hw.mlir:18258:37
    .p0_rd_en   (_T_707),	// matmul/matmul-hw.mlir:18686:13
    .p1_wr_en   (_T_711),	// matmul/matmul-hw.mlir:18673:13
    .p1_wr_data (_T_710),	// matmul/matmul-hw.mlir:18674:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2320)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3424 (	// matmul/matmul-hw.mlir:18259:37
    .p0_rd_en   (_T_702),	// matmul/matmul-hw.mlir:18716:13
    .p1_wr_en   (_T_706),	// matmul/matmul-hw.mlir:18703:13
    .p1_wr_data (_T_705),	// matmul/matmul-hw.mlir:18704:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2319)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3425 (	// matmul/matmul-hw.mlir:18260:37
    .p0_rd_en   (_T_699),	// matmul/matmul-hw.mlir:18743:13
    .p1_wr_en   (_T_701),	// matmul/matmul-hw.mlir:18733:13
    .p1_wr_data (_T_700),	// matmul/matmul-hw.mlir:18734:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2318)
  );
  assign _T_781 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18261:13
  assign _T_780 = _T_2819 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8815:19, :18262:13
  assign _T_779 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18263:13
  assign _T_778 = _T_2808 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18264:13
  mult mult_inst112 (	// matmul/matmul-hw.mlir:18265:28
    .a      (A_reg_bank112_p0_rd_data),	// matmul/matmul-hw.mlir:12327:33
    .b      (_T_2461),
    .t      (_T_2808),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst112_result)
  );
  assign _T_777 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18266:13
  assign a_i_k_0_i_j_7 = A_reg_bank112_p0_rd_data;	// matmul/matmul-hw.mlir:12327:33, :18268:5
  //PROBE: a_i_k_0_i_j_7	// matmul/matmul-hw.mlir:18269:5
  assign b_i_k_0_i_j_7 = _T_2461;	// matmul/matmul-hw.mlir:18271:5
  //PROBE: b_i_k_0_i_j_7	// matmul/matmul-hw.mlir:18272:5
  assign c_prev_i_k_0_i_j_7 = C_reg_bank0_p0_rd_data_2334;	// matmul/matmul-hw.mlir:18244:36, :18274:5
  //PROBE: c_prev_i_k_0_i_j_7	// matmul/matmul-hw.mlir:18275:5
  assign tk_i_k_0_i_j_7 = _T_2786;	// matmul/matmul-hw.mlir:18277:5
  //PROBE: tk_i_k_0_i_j_7	// matmul/matmul-hw.mlir:18278:5
  wire [31:0] _T_3426 = mult_inst112_result + C_reg_bank0_p0_rd_data_2334;	// matmul/matmul-hw.mlir:18244:36, :18265:28, :18279:13
  assign c_i_k_0_i_j_7 = _T_3426;	// matmul/matmul-hw.mlir:18281:5
  //PROBE: c_i_k_0_i_j_7	// matmul/matmul-hw.mlir:18282:5
  assign _T_776 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18283:13
  assign _T_775 = _T_2830 ? _T_3426 : 32'bx;	// matmul/matmul-hw.mlir:8810:19, :18284:13
  localparam [3:0] _T_3428 = 4'h0;	// matmul/matmul-hw.mlir:18287:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18288:5
    if (rst)	// matmul/matmul-hw.mlir:18288:5
      i_k_next_3427 <= _T_3428;	// matmul/matmul-hw.mlir:18291:7
    else	// matmul/matmul-hw.mlir:18288:5
      i_k_next_3427 <= i_j_next_3407;	// matmul/matmul-hw.mlir:18169:13, :18289:7
  end // always @(posedge)
  assign _T_774 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18293:13
  assign _T_773 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18294:13
  mult mult_inst113 (	// matmul/matmul-hw.mlir:18295:28
    .a      (A_reg_bank113_p0_rd_data),	// matmul/matmul-hw.mlir:12328:33
    .b      (_T_2477),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst113_result)
  );
  assign _T_772 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18296:13
  assign a_i_k_1_i_j_7 = A_reg_bank113_p0_rd_data;	// matmul/matmul-hw.mlir:12328:33, :18298:5
  //PROBE: a_i_k_1_i_j_7	// matmul/matmul-hw.mlir:18299:5
  assign b_i_k_1_i_j_7 = _T_2477;	// matmul/matmul-hw.mlir:18301:5
  //PROBE: b_i_k_1_i_j_7	// matmul/matmul-hw.mlir:18302:5
  assign c_prev_i_k_1_i_j_7 = C_reg_bank1_p0_rd_data_2333;	// matmul/matmul-hw.mlir:18245:36, :18304:5
  //PROBE: c_prev_i_k_1_i_j_7	// matmul/matmul-hw.mlir:18305:5
  assign tk_i_k_1_i_j_7 = _T_2797;	// matmul/matmul-hw.mlir:18307:5
  //PROBE: tk_i_k_1_i_j_7	// matmul/matmul-hw.mlir:18308:5
  wire [31:0] _T_3429 = mult_inst113_result + C_reg_bank1_p0_rd_data_2333;	// matmul/matmul-hw.mlir:18245:36, :18295:28, :18309:13
  assign c_i_k_1_i_j_7 = _T_3429;	// matmul/matmul-hw.mlir:18311:5
  //PROBE: c_i_k_1_i_j_7	// matmul/matmul-hw.mlir:18312:5
  assign _T_771 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18313:13
  assign _T_770 = _T_2841 ? _T_3429 : 32'bx;	// matmul/matmul-hw.mlir:8805:19, :18314:13
  localparam [3:0] _T_3431 = 4'h0;	// matmul/matmul-hw.mlir:18317:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18318:5
    if (rst)	// matmul/matmul-hw.mlir:18318:5
      i_k_next_3430 <= _T_3431;	// matmul/matmul-hw.mlir:18321:7
    else	// matmul/matmul-hw.mlir:18318:5
      i_k_next_3430 <= i_k_next_3427;	// matmul/matmul-hw.mlir:18286:13, :18319:7
  end // always @(posedge)
  assign _T_769 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18323:13
  assign _T_768 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18324:13
  mult mult_inst114 (	// matmul/matmul-hw.mlir:18325:28
    .a      (A_reg_bank114_p0_rd_data),	// matmul/matmul-hw.mlir:12329:33
    .b      (_T_2493),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst114_result)
  );
  assign _T_767 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18326:13
  assign a_i_k_2_i_j_7 = A_reg_bank114_p0_rd_data;	// matmul/matmul-hw.mlir:12329:33, :18328:5
  //PROBE: a_i_k_2_i_j_7	// matmul/matmul-hw.mlir:18329:5
  assign b_i_k_2_i_j_7 = _T_2493;	// matmul/matmul-hw.mlir:18331:5
  //PROBE: b_i_k_2_i_j_7	// matmul/matmul-hw.mlir:18332:5
  assign c_prev_i_k_2_i_j_7 = C_reg_bank2_p0_rd_data_2332;	// matmul/matmul-hw.mlir:18246:36, :18334:5
  //PROBE: c_prev_i_k_2_i_j_7	// matmul/matmul-hw.mlir:18335:5
  assign tk_i_k_2_i_j_7 = _T_2808;	// matmul/matmul-hw.mlir:18337:5
  //PROBE: tk_i_k_2_i_j_7	// matmul/matmul-hw.mlir:18338:5
  wire [31:0] _T_3432 = mult_inst114_result + C_reg_bank2_p0_rd_data_2332;	// matmul/matmul-hw.mlir:18246:36, :18325:28, :18339:13
  assign c_i_k_2_i_j_7 = _T_3432;	// matmul/matmul-hw.mlir:18341:5
  //PROBE: c_i_k_2_i_j_7	// matmul/matmul-hw.mlir:18342:5
  assign _T_766 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18343:13
  assign _T_765 = _T_2852 ? _T_3432 : 32'bx;	// matmul/matmul-hw.mlir:8800:19, :18344:13
  localparam [3:0] _T_3434 = 4'h0;	// matmul/matmul-hw.mlir:18347:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18348:5
    if (rst)	// matmul/matmul-hw.mlir:18348:5
      i_k_next_3433 <= _T_3434;	// matmul/matmul-hw.mlir:18351:7
    else	// matmul/matmul-hw.mlir:18348:5
      i_k_next_3433 <= i_k_next_3430;	// matmul/matmul-hw.mlir:18316:13, :18349:7
  end // always @(posedge)
  assign _T_764 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18353:13
  assign _T_763 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18354:13
  mult mult_inst115 (	// matmul/matmul-hw.mlir:18355:28
    .a      (A_reg_bank115_p0_rd_data),	// matmul/matmul-hw.mlir:12330:33
    .b      (_T_2509),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst115_result)
  );
  assign _T_762 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18356:13
  assign a_i_k_3_i_j_7 = A_reg_bank115_p0_rd_data;	// matmul/matmul-hw.mlir:12330:33, :18358:5
  //PROBE: a_i_k_3_i_j_7	// matmul/matmul-hw.mlir:18359:5
  assign b_i_k_3_i_j_7 = _T_2509;	// matmul/matmul-hw.mlir:18361:5
  //PROBE: b_i_k_3_i_j_7	// matmul/matmul-hw.mlir:18362:5
  assign c_prev_i_k_3_i_j_7 = C_reg_bank3_p0_rd_data_2331;	// matmul/matmul-hw.mlir:18247:36, :18364:5
  //PROBE: c_prev_i_k_3_i_j_7	// matmul/matmul-hw.mlir:18365:5
  assign tk_i_k_3_i_j_7 = _T_2819;	// matmul/matmul-hw.mlir:18367:5
  //PROBE: tk_i_k_3_i_j_7	// matmul/matmul-hw.mlir:18368:5
  wire [31:0] _T_3435 = mult_inst115_result + C_reg_bank3_p0_rd_data_2331;	// matmul/matmul-hw.mlir:18247:36, :18355:28, :18369:13
  assign c_i_k_3_i_j_7 = _T_3435;	// matmul/matmul-hw.mlir:18371:5
  //PROBE: c_i_k_3_i_j_7	// matmul/matmul-hw.mlir:18372:5
  assign _T_761 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18373:13
  assign _T_760 = _T_2863 ? _T_3435 : 32'bx;	// matmul/matmul-hw.mlir:8795:19, :18374:13
  localparam [3:0] _T_3437 = 4'h0;	// matmul/matmul-hw.mlir:18377:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18378:5
    if (rst)	// matmul/matmul-hw.mlir:18378:5
      i_k_next_3436 <= _T_3437;	// matmul/matmul-hw.mlir:18381:7
    else	// matmul/matmul-hw.mlir:18378:5
      i_k_next_3436 <= i_k_next_3433;	// matmul/matmul-hw.mlir:18346:13, :18379:7
  end // always @(posedge)
  assign _T_759 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18383:13
  assign _T_758 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18384:13
  mult mult_inst116 (	// matmul/matmul-hw.mlir:18385:28
    .a      (A_reg_bank116_p0_rd_data),	// matmul/matmul-hw.mlir:12331:33
    .b      (_T_2525),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst116_result)
  );
  assign _T_757 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18386:13
  assign a_i_k_4_i_j_7 = A_reg_bank116_p0_rd_data;	// matmul/matmul-hw.mlir:12331:33, :18388:5
  //PROBE: a_i_k_4_i_j_7	// matmul/matmul-hw.mlir:18389:5
  assign b_i_k_4_i_j_7 = _T_2525;	// matmul/matmul-hw.mlir:18391:5
  //PROBE: b_i_k_4_i_j_7	// matmul/matmul-hw.mlir:18392:5
  assign c_prev_i_k_4_i_j_7 = C_reg_bank4_p0_rd_data_2330;	// matmul/matmul-hw.mlir:18248:36, :18394:5
  //PROBE: c_prev_i_k_4_i_j_7	// matmul/matmul-hw.mlir:18395:5
  assign tk_i_k_4_i_j_7 = _T_2830;	// matmul/matmul-hw.mlir:18397:5
  //PROBE: tk_i_k_4_i_j_7	// matmul/matmul-hw.mlir:18398:5
  wire [31:0] _T_3438 = mult_inst116_result + C_reg_bank4_p0_rd_data_2330;	// matmul/matmul-hw.mlir:18248:36, :18385:28, :18399:13
  assign c_i_k_4_i_j_7 = _T_3438;	// matmul/matmul-hw.mlir:18401:5
  //PROBE: c_i_k_4_i_j_7	// matmul/matmul-hw.mlir:18402:5
  assign _T_756 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18403:13
  assign _T_755 = _T_2874 ? _T_3438 : 32'bx;	// matmul/matmul-hw.mlir:8790:19, :18404:13
  localparam [3:0] _T_3440 = 4'h0;	// matmul/matmul-hw.mlir:18407:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18408:5
    if (rst)	// matmul/matmul-hw.mlir:18408:5
      i_k_next_3439 <= _T_3440;	// matmul/matmul-hw.mlir:18411:7
    else	// matmul/matmul-hw.mlir:18408:5
      i_k_next_3439 <= i_k_next_3436;	// matmul/matmul-hw.mlir:18376:13, :18409:7
  end // always @(posedge)
  assign _T_754 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18413:13
  assign _T_753 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18414:13
  mult mult_inst117 (	// matmul/matmul-hw.mlir:18415:28
    .a      (A_reg_bank117_p0_rd_data),	// matmul/matmul-hw.mlir:12332:33
    .b      (_T_2541),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst117_result)
  );
  assign _T_752 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18416:13
  assign a_i_k_5_i_j_7 = A_reg_bank117_p0_rd_data;	// matmul/matmul-hw.mlir:12332:33, :18418:5
  //PROBE: a_i_k_5_i_j_7	// matmul/matmul-hw.mlir:18419:5
  assign b_i_k_5_i_j_7 = _T_2541;	// matmul/matmul-hw.mlir:18421:5
  //PROBE: b_i_k_5_i_j_7	// matmul/matmul-hw.mlir:18422:5
  assign c_prev_i_k_5_i_j_7 = C_reg_bank5_p0_rd_data_2329;	// matmul/matmul-hw.mlir:18249:36, :18424:5
  //PROBE: c_prev_i_k_5_i_j_7	// matmul/matmul-hw.mlir:18425:5
  assign tk_i_k_5_i_j_7 = _T_2841;	// matmul/matmul-hw.mlir:18427:5
  //PROBE: tk_i_k_5_i_j_7	// matmul/matmul-hw.mlir:18428:5
  wire [31:0] _T_3441 = mult_inst117_result + C_reg_bank5_p0_rd_data_2329;	// matmul/matmul-hw.mlir:18249:36, :18415:28, :18429:13
  assign c_i_k_5_i_j_7 = _T_3441;	// matmul/matmul-hw.mlir:18431:5
  //PROBE: c_i_k_5_i_j_7	// matmul/matmul-hw.mlir:18432:5
  assign _T_751 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18433:13
  assign _T_750 = _T_2885 ? _T_3441 : 32'bx;	// matmul/matmul-hw.mlir:8785:19, :18434:13
  localparam [3:0] _T_3443 = 4'h0;	// matmul/matmul-hw.mlir:18437:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18438:5
    if (rst)	// matmul/matmul-hw.mlir:18438:5
      i_k_next_3442 <= _T_3443;	// matmul/matmul-hw.mlir:18441:7
    else	// matmul/matmul-hw.mlir:18438:5
      i_k_next_3442 <= i_k_next_3439;	// matmul/matmul-hw.mlir:18406:13, :18439:7
  end // always @(posedge)
  assign _T_749 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18443:13
  assign _T_748 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18444:13
  mult mult_inst118 (	// matmul/matmul-hw.mlir:18445:28
    .a      (A_reg_bank118_p0_rd_data),	// matmul/matmul-hw.mlir:12333:33
    .b      (_T_2557),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst118_result)
  );
  assign _T_747 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18446:13
  assign a_i_k_6_i_j_7 = A_reg_bank118_p0_rd_data;	// matmul/matmul-hw.mlir:12333:33, :18448:5
  //PROBE: a_i_k_6_i_j_7	// matmul/matmul-hw.mlir:18449:5
  assign b_i_k_6_i_j_7 = _T_2557;	// matmul/matmul-hw.mlir:18451:5
  //PROBE: b_i_k_6_i_j_7	// matmul/matmul-hw.mlir:18452:5
  assign c_prev_i_k_6_i_j_7 = C_reg_bank6_p0_rd_data_2328;	// matmul/matmul-hw.mlir:18250:36, :18454:5
  //PROBE: c_prev_i_k_6_i_j_7	// matmul/matmul-hw.mlir:18455:5
  assign tk_i_k_6_i_j_7 = _T_2852;	// matmul/matmul-hw.mlir:18457:5
  //PROBE: tk_i_k_6_i_j_7	// matmul/matmul-hw.mlir:18458:5
  wire [31:0] _T_3444 = mult_inst118_result + C_reg_bank6_p0_rd_data_2328;	// matmul/matmul-hw.mlir:18250:36, :18445:28, :18459:13
  assign c_i_k_6_i_j_7 = _T_3444;	// matmul/matmul-hw.mlir:18461:5
  //PROBE: c_i_k_6_i_j_7	// matmul/matmul-hw.mlir:18462:5
  assign _T_746 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18463:13
  assign _T_745 = _T_2892 ? _T_3444 : 32'bx;	// matmul/matmul-hw.mlir:8780:19, :18464:13
  localparam [3:0] _T_3446 = 4'h0;	// matmul/matmul-hw.mlir:18467:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18468:5
    if (rst)	// matmul/matmul-hw.mlir:18468:5
      i_k_next_3445 <= _T_3446;	// matmul/matmul-hw.mlir:18471:7
    else	// matmul/matmul-hw.mlir:18468:5
      i_k_next_3445 <= i_k_next_3442;	// matmul/matmul-hw.mlir:18436:13, :18469:7
  end // always @(posedge)
  assign _T_744 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18473:13
  assign _T_743 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18474:13
  mult mult_inst119 (	// matmul/matmul-hw.mlir:18475:28
    .a      (A_reg_bank119_p0_rd_data),	// matmul/matmul-hw.mlir:12334:33
    .b      (_T_2573),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst119_result)
  );
  assign _T_742 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18476:13
  assign a_i_k_7_i_j_7 = A_reg_bank119_p0_rd_data;	// matmul/matmul-hw.mlir:12334:33, :18478:5
  //PROBE: a_i_k_7_i_j_7	// matmul/matmul-hw.mlir:18479:5
  assign b_i_k_7_i_j_7 = _T_2573;	// matmul/matmul-hw.mlir:18481:5
  //PROBE: b_i_k_7_i_j_7	// matmul/matmul-hw.mlir:18482:5
  assign c_prev_i_k_7_i_j_7 = C_reg_bank7_p0_rd_data_2327;	// matmul/matmul-hw.mlir:18251:36, :18484:5
  //PROBE: c_prev_i_k_7_i_j_7	// matmul/matmul-hw.mlir:18485:5
  assign tk_i_k_7_i_j_7 = _T_2863;	// matmul/matmul-hw.mlir:18487:5
  //PROBE: tk_i_k_7_i_j_7	// matmul/matmul-hw.mlir:18488:5
  wire [31:0] _T_3447 = mult_inst119_result + C_reg_bank7_p0_rd_data_2327;	// matmul/matmul-hw.mlir:18251:36, :18475:28, :18489:13
  assign c_i_k_7_i_j_7 = _T_3447;	// matmul/matmul-hw.mlir:18491:5
  //PROBE: c_i_k_7_i_j_7	// matmul/matmul-hw.mlir:18492:5
  assign _T_741 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18493:13
  assign _T_740 = _T_2897 ? _T_3447 : 32'bx;	// matmul/matmul-hw.mlir:8775:19, :18494:13
  localparam [3:0] _T_3449 = 4'h0;	// matmul/matmul-hw.mlir:18497:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18498:5
    if (rst)	// matmul/matmul-hw.mlir:18498:5
      i_k_next_3448 <= _T_3449;	// matmul/matmul-hw.mlir:18501:7
    else	// matmul/matmul-hw.mlir:18498:5
      i_k_next_3448 <= i_k_next_3445;	// matmul/matmul-hw.mlir:18466:13, :18499:7
  end // always @(posedge)
  assign _T_739 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18503:13
  assign _T_738 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18504:13
  mult mult_inst120 (	// matmul/matmul-hw.mlir:18505:28
    .a      (A_reg_bank120_p0_rd_data),	// matmul/matmul-hw.mlir:12335:33
    .b      (_T_2589),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst120_result)
  );
  assign _T_737 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18506:13
  assign a_i_k_8_i_j_7 = A_reg_bank120_p0_rd_data;	// matmul/matmul-hw.mlir:12335:33, :18508:5
  //PROBE: a_i_k_8_i_j_7	// matmul/matmul-hw.mlir:18509:5
  assign b_i_k_8_i_j_7 = _T_2589;	// matmul/matmul-hw.mlir:18511:5
  //PROBE: b_i_k_8_i_j_7	// matmul/matmul-hw.mlir:18512:5
  assign c_prev_i_k_8_i_j_7 = C_reg_bank8_p0_rd_data_2326;	// matmul/matmul-hw.mlir:18252:36, :18514:5
  //PROBE: c_prev_i_k_8_i_j_7	// matmul/matmul-hw.mlir:18515:5
  assign tk_i_k_8_i_j_7 = _T_2874;	// matmul/matmul-hw.mlir:18517:5
  //PROBE: tk_i_k_8_i_j_7	// matmul/matmul-hw.mlir:18518:5
  wire [31:0] _T_3450 = mult_inst120_result + C_reg_bank8_p0_rd_data_2326;	// matmul/matmul-hw.mlir:18252:36, :18505:28, :18519:13
  assign c_i_k_8_i_j_7 = _T_3450;	// matmul/matmul-hw.mlir:18521:5
  //PROBE: c_i_k_8_i_j_7	// matmul/matmul-hw.mlir:18522:5
  assign _T_736 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18523:13
  assign _T_735 = _T_2902 ? _T_3450 : 32'bx;	// matmul/matmul-hw.mlir:8770:19, :18524:13
  localparam [3:0] _T_3452 = 4'h0;	// matmul/matmul-hw.mlir:18527:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18528:5
    if (rst)	// matmul/matmul-hw.mlir:18528:5
      i_k_next_3451 <= _T_3452;	// matmul/matmul-hw.mlir:18531:7
    else	// matmul/matmul-hw.mlir:18528:5
      i_k_next_3451 <= i_k_next_3448;	// matmul/matmul-hw.mlir:18496:13, :18529:7
  end // always @(posedge)
  assign _T_734 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18533:13
  assign _T_733 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18534:13
  mult mult_inst121 (	// matmul/matmul-hw.mlir:18535:28
    .a      (A_reg_bank121_p0_rd_data),	// matmul/matmul-hw.mlir:12336:33
    .b      (_T_2605),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst121_result)
  );
  assign _T_732 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18536:13
  assign a_i_k_9_i_j_7 = A_reg_bank121_p0_rd_data;	// matmul/matmul-hw.mlir:12336:33, :18538:5
  //PROBE: a_i_k_9_i_j_7	// matmul/matmul-hw.mlir:18539:5
  assign b_i_k_9_i_j_7 = _T_2605;	// matmul/matmul-hw.mlir:18541:5
  //PROBE: b_i_k_9_i_j_7	// matmul/matmul-hw.mlir:18542:5
  assign c_prev_i_k_9_i_j_7 = C_reg_bank9_p0_rd_data_2325;	// matmul/matmul-hw.mlir:18253:36, :18544:5
  //PROBE: c_prev_i_k_9_i_j_7	// matmul/matmul-hw.mlir:18545:5
  assign tk_i_k_9_i_j_7 = _T_2885;	// matmul/matmul-hw.mlir:18547:5
  //PROBE: tk_i_k_9_i_j_7	// matmul/matmul-hw.mlir:18548:5
  wire [31:0] _T_3453 = mult_inst121_result + C_reg_bank9_p0_rd_data_2325;	// matmul/matmul-hw.mlir:18253:36, :18535:28, :18549:13
  assign c_i_k_9_i_j_7 = _T_3453;	// matmul/matmul-hw.mlir:18551:5
  //PROBE: c_i_k_9_i_j_7	// matmul/matmul-hw.mlir:18552:5
  assign _T_731 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18553:13
  assign _T_730 = _T_2907 ? _T_3453 : 32'bx;	// matmul/matmul-hw.mlir:8765:19, :18554:13
  localparam [3:0] _T_3455 = 4'h0;	// matmul/matmul-hw.mlir:18557:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18558:5
    if (rst)	// matmul/matmul-hw.mlir:18558:5
      i_k_next_3454 <= _T_3455;	// matmul/matmul-hw.mlir:18561:7
    else	// matmul/matmul-hw.mlir:18558:5
      i_k_next_3454 <= i_k_next_3451;	// matmul/matmul-hw.mlir:18526:13, :18559:7
  end // always @(posedge)
  assign _T_729 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18563:13
  assign _T_728 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18564:13
  mult mult_inst122 (	// matmul/matmul-hw.mlir:18565:28
    .a      (A_reg_bank122_p0_rd_data),	// matmul/matmul-hw.mlir:12337:33
    .b      (_T_2621),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst122_result)
  );
  assign _T_727 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18566:13
  assign a_i_k_10_i_j_7 = A_reg_bank122_p0_rd_data;	// matmul/matmul-hw.mlir:12337:33, :18568:5
  //PROBE: a_i_k_10_i_j_7	// matmul/matmul-hw.mlir:18569:5
  assign b_i_k_10_i_j_7 = _T_2621;	// matmul/matmul-hw.mlir:18571:5
  //PROBE: b_i_k_10_i_j_7	// matmul/matmul-hw.mlir:18572:5
  assign c_prev_i_k_10_i_j_7 = C_reg_bank10_p0_rd_data_2324;	// matmul/matmul-hw.mlir:18254:37, :18574:5
  //PROBE: c_prev_i_k_10_i_j_7	// matmul/matmul-hw.mlir:18575:5
  assign tk_i_k_10_i_j_7 = _T_2892;	// matmul/matmul-hw.mlir:18577:5
  //PROBE: tk_i_k_10_i_j_7	// matmul/matmul-hw.mlir:18578:5
  wire [31:0] _T_3456 = mult_inst122_result + C_reg_bank10_p0_rd_data_2324;	// matmul/matmul-hw.mlir:18254:37, :18565:28, :18579:13
  assign c_i_k_10_i_j_7 = _T_3456;	// matmul/matmul-hw.mlir:18581:5
  //PROBE: c_i_k_10_i_j_7	// matmul/matmul-hw.mlir:18582:5
  assign _T_726 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18583:13
  assign _T_725 = _T_2912 ? _T_3456 : 32'bx;	// matmul/matmul-hw.mlir:8760:19, :18584:13
  localparam [3:0] _T_3458 = 4'h0;	// matmul/matmul-hw.mlir:18587:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18588:5
    if (rst)	// matmul/matmul-hw.mlir:18588:5
      i_k_next_3457 <= _T_3458;	// matmul/matmul-hw.mlir:18591:7
    else	// matmul/matmul-hw.mlir:18588:5
      i_k_next_3457 <= i_k_next_3454;	// matmul/matmul-hw.mlir:18556:13, :18589:7
  end // always @(posedge)
  assign _T_724 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18593:13
  assign _T_723 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18594:13
  mult mult_inst123 (	// matmul/matmul-hw.mlir:18595:28
    .a      (A_reg_bank123_p0_rd_data),	// matmul/matmul-hw.mlir:12338:33
    .b      (_T_2637),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst123_result)
  );
  assign _T_722 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18596:13
  assign a_i_k_11_i_j_7 = A_reg_bank123_p0_rd_data;	// matmul/matmul-hw.mlir:12338:33, :18598:5
  //PROBE: a_i_k_11_i_j_7	// matmul/matmul-hw.mlir:18599:5
  assign b_i_k_11_i_j_7 = _T_2637;	// matmul/matmul-hw.mlir:18601:5
  //PROBE: b_i_k_11_i_j_7	// matmul/matmul-hw.mlir:18602:5
  assign c_prev_i_k_11_i_j_7 = C_reg_bank11_p0_rd_data_2323;	// matmul/matmul-hw.mlir:18255:37, :18604:5
  //PROBE: c_prev_i_k_11_i_j_7	// matmul/matmul-hw.mlir:18605:5
  assign tk_i_k_11_i_j_7 = _T_2897;	// matmul/matmul-hw.mlir:18607:5
  //PROBE: tk_i_k_11_i_j_7	// matmul/matmul-hw.mlir:18608:5
  wire [31:0] _T_3459 = mult_inst123_result + C_reg_bank11_p0_rd_data_2323;	// matmul/matmul-hw.mlir:18255:37, :18595:28, :18609:13
  assign c_i_k_11_i_j_7 = _T_3459;	// matmul/matmul-hw.mlir:18611:5
  //PROBE: c_i_k_11_i_j_7	// matmul/matmul-hw.mlir:18612:5
  assign _T_721 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18613:13
  assign _T_720 = _T_2917 ? _T_3459 : 32'bx;	// matmul/matmul-hw.mlir:8755:19, :18614:13
  localparam [3:0] _T_3461 = 4'h0;	// matmul/matmul-hw.mlir:18617:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18618:5
    if (rst)	// matmul/matmul-hw.mlir:18618:5
      i_k_next_3460 <= _T_3461;	// matmul/matmul-hw.mlir:18621:7
    else	// matmul/matmul-hw.mlir:18618:5
      i_k_next_3460 <= i_k_next_3457;	// matmul/matmul-hw.mlir:18586:13, :18619:7
  end // always @(posedge)
  assign _T_719 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18623:13
  assign _T_718 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18624:13
  mult mult_inst124 (	// matmul/matmul-hw.mlir:18625:28
    .a      (A_reg_bank124_p0_rd_data),	// matmul/matmul-hw.mlir:12339:33
    .b      (_T_2653),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst124_result)
  );
  assign _T_717 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18626:13
  assign a_i_k_12_i_j_7 = A_reg_bank124_p0_rd_data;	// matmul/matmul-hw.mlir:12339:33, :18628:5
  //PROBE: a_i_k_12_i_j_7	// matmul/matmul-hw.mlir:18629:5
  assign b_i_k_12_i_j_7 = _T_2653;	// matmul/matmul-hw.mlir:18631:5
  //PROBE: b_i_k_12_i_j_7	// matmul/matmul-hw.mlir:18632:5
  assign c_prev_i_k_12_i_j_7 = C_reg_bank12_p0_rd_data_2322;	// matmul/matmul-hw.mlir:18256:37, :18634:5
  //PROBE: c_prev_i_k_12_i_j_7	// matmul/matmul-hw.mlir:18635:5
  assign tk_i_k_12_i_j_7 = _T_2902;	// matmul/matmul-hw.mlir:18637:5
  //PROBE: tk_i_k_12_i_j_7	// matmul/matmul-hw.mlir:18638:5
  wire [31:0] _T_3462 = mult_inst124_result + C_reg_bank12_p0_rd_data_2322;	// matmul/matmul-hw.mlir:18256:37, :18625:28, :18639:13
  assign c_i_k_12_i_j_7 = _T_3462;	// matmul/matmul-hw.mlir:18641:5
  //PROBE: c_i_k_12_i_j_7	// matmul/matmul-hw.mlir:18642:5
  assign _T_716 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18643:13
  assign _T_715 = _T_2922 ? _T_3462 : 32'bx;	// matmul/matmul-hw.mlir:8750:19, :18644:13
  localparam [3:0] _T_3464 = 4'h0;	// matmul/matmul-hw.mlir:18647:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18648:5
    if (rst)	// matmul/matmul-hw.mlir:18648:5
      i_k_next_3463 <= _T_3464;	// matmul/matmul-hw.mlir:18651:7
    else	// matmul/matmul-hw.mlir:18648:5
      i_k_next_3463 <= i_k_next_3460;	// matmul/matmul-hw.mlir:18616:13, :18649:7
  end // always @(posedge)
  assign _T_714 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18653:13
  assign _T_713 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18654:13
  mult mult_inst125 (	// matmul/matmul-hw.mlir:18655:28
    .a      (A_reg_bank125_p0_rd_data),	// matmul/matmul-hw.mlir:12340:33
    .b      (_T_2669),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst125_result)
  );
  assign _T_712 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18656:13
  assign a_i_k_13_i_j_7 = A_reg_bank125_p0_rd_data;	// matmul/matmul-hw.mlir:12340:33, :18658:5
  //PROBE: a_i_k_13_i_j_7	// matmul/matmul-hw.mlir:18659:5
  assign b_i_k_13_i_j_7 = _T_2669;	// matmul/matmul-hw.mlir:18661:5
  //PROBE: b_i_k_13_i_j_7	// matmul/matmul-hw.mlir:18662:5
  assign c_prev_i_k_13_i_j_7 = C_reg_bank13_p0_rd_data_2321;	// matmul/matmul-hw.mlir:18257:37, :18664:5
  //PROBE: c_prev_i_k_13_i_j_7	// matmul/matmul-hw.mlir:18665:5
  assign tk_i_k_13_i_j_7 = _T_2907;	// matmul/matmul-hw.mlir:18667:5
  //PROBE: tk_i_k_13_i_j_7	// matmul/matmul-hw.mlir:18668:5
  wire [31:0] _T_3465 = mult_inst125_result + C_reg_bank13_p0_rd_data_2321;	// matmul/matmul-hw.mlir:18257:37, :18655:28, :18669:13
  assign c_i_k_13_i_j_7 = _T_3465;	// matmul/matmul-hw.mlir:18671:5
  //PROBE: c_i_k_13_i_j_7	// matmul/matmul-hw.mlir:18672:5
  assign _T_711 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18673:13
  assign _T_710 = _T_2927 ? _T_3465 : 32'bx;	// matmul/matmul-hw.mlir:8745:19, :18674:13
  localparam [3:0] _T_3467 = 4'h0;	// matmul/matmul-hw.mlir:18677:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18678:5
    if (rst)	// matmul/matmul-hw.mlir:18678:5
      i_k_next_3466 <= _T_3467;	// matmul/matmul-hw.mlir:18681:7
    else	// matmul/matmul-hw.mlir:18678:5
      i_k_next_3466 <= i_k_next_3463;	// matmul/matmul-hw.mlir:18646:13, :18679:7
  end // always @(posedge)
  assign _T_709 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18683:13
  assign _T_708 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18684:13
  mult mult_inst126 (	// matmul/matmul-hw.mlir:18685:28
    .a      (A_reg_bank126_p0_rd_data),	// matmul/matmul-hw.mlir:12341:33
    .b      (_T_2685),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst126_result)
  );
  assign _T_707 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18686:13
  assign a_i_k_14_i_j_7 = A_reg_bank126_p0_rd_data;	// matmul/matmul-hw.mlir:12341:33, :18688:5
  //PROBE: a_i_k_14_i_j_7	// matmul/matmul-hw.mlir:18689:5
  assign b_i_k_14_i_j_7 = _T_2685;	// matmul/matmul-hw.mlir:18691:5
  //PROBE: b_i_k_14_i_j_7	// matmul/matmul-hw.mlir:18692:5
  assign c_prev_i_k_14_i_j_7 = C_reg_bank14_p0_rd_data_2320;	// matmul/matmul-hw.mlir:18258:37, :18694:5
  //PROBE: c_prev_i_k_14_i_j_7	// matmul/matmul-hw.mlir:18695:5
  assign tk_i_k_14_i_j_7 = _T_2912;	// matmul/matmul-hw.mlir:18697:5
  //PROBE: tk_i_k_14_i_j_7	// matmul/matmul-hw.mlir:18698:5
  wire [31:0] _T_3468 = mult_inst126_result + C_reg_bank14_p0_rd_data_2320;	// matmul/matmul-hw.mlir:18258:37, :18685:28, :18699:13
  assign c_i_k_14_i_j_7 = _T_3468;	// matmul/matmul-hw.mlir:18701:5
  //PROBE: c_i_k_14_i_j_7	// matmul/matmul-hw.mlir:18702:5
  assign _T_706 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18703:13
  assign _T_705 = _T_2932 ? _T_3468 : 32'bx;	// matmul/matmul-hw.mlir:8740:19, :18704:13
  localparam [3:0] _T_3470 = 4'h0;	// matmul/matmul-hw.mlir:18707:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18708:5
    if (rst)	// matmul/matmul-hw.mlir:18708:5
      i_k_next_3469 <= _T_3470;	// matmul/matmul-hw.mlir:18711:7
    else	// matmul/matmul-hw.mlir:18708:5
      i_k_next_3469 <= i_k_next_3466;	// matmul/matmul-hw.mlir:18676:13, :18709:7
  end // always @(posedge)
  assign _T_704 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18713:13
  assign _T_703 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18714:13
  mult mult_inst127 (	// matmul/matmul-hw.mlir:18715:28
    .a      (A_reg_bank127_p0_rd_data),	// matmul/matmul-hw.mlir:12342:33
    .b      (_T_2701),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst127_result)
  );
  assign _T_702 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18716:13
  assign a_i_k_15_i_j_7 = A_reg_bank127_p0_rd_data;	// matmul/matmul-hw.mlir:12342:33, :18718:5
  //PROBE: a_i_k_15_i_j_7	// matmul/matmul-hw.mlir:18719:5
  assign b_i_k_15_i_j_7 = _T_2701;	// matmul/matmul-hw.mlir:18721:5
  //PROBE: b_i_k_15_i_j_7	// matmul/matmul-hw.mlir:18722:5
  assign c_prev_i_k_15_i_j_7 = C_reg_bank15_p0_rd_data_2319;	// matmul/matmul-hw.mlir:18259:37, :18724:5
  //PROBE: c_prev_i_k_15_i_j_7	// matmul/matmul-hw.mlir:18725:5
  assign tk_i_k_15_i_j_7 = _T_2917;	// matmul/matmul-hw.mlir:18727:5
  //PROBE: tk_i_k_15_i_j_7	// matmul/matmul-hw.mlir:18728:5
  wire [31:0] _T_3471 = mult_inst127_result + C_reg_bank15_p0_rd_data_2319;	// matmul/matmul-hw.mlir:18259:37, :18715:28, :18729:13
  assign c_i_k_15_i_j_7 = _T_3471;	// matmul/matmul-hw.mlir:18731:5
  //PROBE: c_i_k_15_i_j_7	// matmul/matmul-hw.mlir:18732:5
  assign _T_701 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18733:13
  assign _T_700 = _T_2937 ? _T_3471 : 32'bx;	// matmul/matmul-hw.mlir:8735:19, :18734:13
  localparam [3:0] _T_3473 = 4'h0;	// matmul/matmul-hw.mlir:18737:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18738:5
    if (rst)	// matmul/matmul-hw.mlir:18738:5
      i_k_next_3472 <= _T_3473;	// matmul/matmul-hw.mlir:18741:7
    else	// matmul/matmul-hw.mlir:18738:5
      i_k_next_3472 <= i_k_next_3469;	// matmul/matmul-hw.mlir:18706:13, :18739:7
  end // always @(posedge)
  assign _T_699 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18743:13
  wire [3:0][3:0] _T_3475 = i_delayed_3474;	// matmul/matmul-hw.mlir:18745:13
  wire [3:0][3:0] _T_3476 = {_T_3475[2'h0+:3], {{i_k_next_3472}}};	// matmul/matmul-hw.mlir:18736:13, :18746:19, :18747:13, :18748:13, :18749:13
  wire [3:0][3:0] _T_3477 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:18750:19, :18751:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18752:5
    if (rst)	// matmul/matmul-hw.mlir:18752:5
      i_delayed_3474 <= _T_3477;	// matmul/matmul-hw.mlir:18755:7
    else	// matmul/matmul-hw.mlir:18752:5
      i_delayed_3474 <= _T_3476;	// matmul/matmul-hw.mlir:18753:7
  end // always @(posedge)
  assign _T_698 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18759:13
  assign _T_697 = _T_2942 ? i_delayed_3474[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8732:18, :18745:13, :18757:20, :18758:13, :18760:13
  assign _T_696 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18761:13
  assign _T_695 = _T_2942 ? C_reg_bank16_p0_rd_data_2318 : 32'bx;	// matmul/matmul-hw.mlir:8730:19, :18260:37, :18762:13
  localparam [3:0] _T_3479 = 4'h0;	// matmul/matmul-hw.mlir:18765:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18766:5
    if (rst)	// matmul/matmul-hw.mlir:18766:5
      i_j_next_3478 <= _T_3479;	// matmul/matmul-hw.mlir:18769:7
    else	// matmul/matmul-hw.mlir:18766:5
      i_j_next_3478 <= i_j_next_3407;	// matmul/matmul-hw.mlir:18169:13, :18767:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3480 (	// matmul/matmul-hw.mlir:18839:36
    .p0_rd_en   (_T_690),	// matmul/matmul-hw.mlir:18861:13
    .p1_wr_en   (_T_694),	// matmul/matmul-hw.mlir:18856:13
    .p1_wr_data (_T_693),	// matmul/matmul-hw.mlir:18857:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2317)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3481 (	// matmul/matmul-hw.mlir:18840:36
    .p0_rd_en   (_T_685),	// matmul/matmul-hw.mlir:18891:13
    .p1_wr_en   (_T_689),	// matmul/matmul-hw.mlir:18878:13
    .p1_wr_data (_T_688),	// matmul/matmul-hw.mlir:18879:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2316)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3482 (	// matmul/matmul-hw.mlir:18841:36
    .p0_rd_en   (_T_680),	// matmul/matmul-hw.mlir:18921:13
    .p1_wr_en   (_T_684),	// matmul/matmul-hw.mlir:18908:13
    .p1_wr_data (_T_683),	// matmul/matmul-hw.mlir:18909:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2315)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3483 (	// matmul/matmul-hw.mlir:18842:36
    .p0_rd_en   (_T_675),	// matmul/matmul-hw.mlir:18951:13
    .p1_wr_en   (_T_679),	// matmul/matmul-hw.mlir:18938:13
    .p1_wr_data (_T_678),	// matmul/matmul-hw.mlir:18939:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2314)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3484 (	// matmul/matmul-hw.mlir:18843:36
    .p0_rd_en   (_T_670),	// matmul/matmul-hw.mlir:18981:13
    .p1_wr_en   (_T_674),	// matmul/matmul-hw.mlir:18968:13
    .p1_wr_data (_T_673),	// matmul/matmul-hw.mlir:18969:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2313)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3485 (	// matmul/matmul-hw.mlir:18844:36
    .p0_rd_en   (_T_665),	// matmul/matmul-hw.mlir:19011:13
    .p1_wr_en   (_T_669),	// matmul/matmul-hw.mlir:18998:13
    .p1_wr_data (_T_668),	// matmul/matmul-hw.mlir:18999:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2312)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3486 (	// matmul/matmul-hw.mlir:18845:36
    .p0_rd_en   (_T_660),	// matmul/matmul-hw.mlir:19041:13
    .p1_wr_en   (_T_664),	// matmul/matmul-hw.mlir:19028:13
    .p1_wr_data (_T_663),	// matmul/matmul-hw.mlir:19029:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2311)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3487 (	// matmul/matmul-hw.mlir:18846:36
    .p0_rd_en   (_T_655),	// matmul/matmul-hw.mlir:19071:13
    .p1_wr_en   (_T_659),	// matmul/matmul-hw.mlir:19058:13
    .p1_wr_data (_T_658),	// matmul/matmul-hw.mlir:19059:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2310)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3488 (	// matmul/matmul-hw.mlir:18847:36
    .p0_rd_en   (_T_650),	// matmul/matmul-hw.mlir:19101:13
    .p1_wr_en   (_T_654),	// matmul/matmul-hw.mlir:19088:13
    .p1_wr_data (_T_653),	// matmul/matmul-hw.mlir:19089:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2309)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3489 (	// matmul/matmul-hw.mlir:18848:36
    .p0_rd_en   (_T_645),	// matmul/matmul-hw.mlir:19131:13
    .p1_wr_en   (_T_649),	// matmul/matmul-hw.mlir:19118:13
    .p1_wr_data (_T_648),	// matmul/matmul-hw.mlir:19119:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2308)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3490 (	// matmul/matmul-hw.mlir:18849:37
    .p0_rd_en   (_T_640),	// matmul/matmul-hw.mlir:19161:13
    .p1_wr_en   (_T_644),	// matmul/matmul-hw.mlir:19148:13
    .p1_wr_data (_T_643),	// matmul/matmul-hw.mlir:19149:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2307)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3491 (	// matmul/matmul-hw.mlir:18850:37
    .p0_rd_en   (_T_635),	// matmul/matmul-hw.mlir:19191:13
    .p1_wr_en   (_T_639),	// matmul/matmul-hw.mlir:19178:13
    .p1_wr_data (_T_638),	// matmul/matmul-hw.mlir:19179:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2306)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3492 (	// matmul/matmul-hw.mlir:18851:37
    .p0_rd_en   (_T_630),	// matmul/matmul-hw.mlir:19221:13
    .p1_wr_en   (_T_634),	// matmul/matmul-hw.mlir:19208:13
    .p1_wr_data (_T_633),	// matmul/matmul-hw.mlir:19209:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2305)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3493 (	// matmul/matmul-hw.mlir:18852:37
    .p0_rd_en   (_T_625),	// matmul/matmul-hw.mlir:19251:13
    .p1_wr_en   (_T_629),	// matmul/matmul-hw.mlir:19238:13
    .p1_wr_data (_T_628),	// matmul/matmul-hw.mlir:19239:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2304)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3494 (	// matmul/matmul-hw.mlir:18853:37
    .p0_rd_en   (_T_620),	// matmul/matmul-hw.mlir:19281:13
    .p1_wr_en   (_T_624),	// matmul/matmul-hw.mlir:19268:13
    .p1_wr_data (_T_623),	// matmul/matmul-hw.mlir:19269:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2303)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3495 (	// matmul/matmul-hw.mlir:18854:37
    .p0_rd_en   (_T_615),	// matmul/matmul-hw.mlir:19311:13
    .p1_wr_en   (_T_619),	// matmul/matmul-hw.mlir:19298:13
    .p1_wr_data (_T_618),	// matmul/matmul-hw.mlir:19299:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2302)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3496 (	// matmul/matmul-hw.mlir:18855:37
    .p0_rd_en   (_T_612),	// matmul/matmul-hw.mlir:19338:13
    .p1_wr_en   (_T_614),	// matmul/matmul-hw.mlir:19328:13
    .p1_wr_data (_T_613),	// matmul/matmul-hw.mlir:19329:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2301)
  );
  assign _T_694 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18856:13
  assign _T_693 = _T_2830 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8728:19, :18857:13
  assign _T_692 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18858:13
  assign _T_691 = _T_2819 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18859:13
  mult mult_inst128 (	// matmul/matmul-hw.mlir:18860:28
    .a      (A_reg_bank128_p0_rd_data),	// matmul/matmul-hw.mlir:12343:33
    .b      (_T_2462),
    .t      (_T_2819),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst128_result)
  );
  assign _T_690 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18861:13
  assign a_i_k_0_i_j_8 = A_reg_bank128_p0_rd_data;	// matmul/matmul-hw.mlir:12343:33, :18863:5
  //PROBE: a_i_k_0_i_j_8	// matmul/matmul-hw.mlir:18864:5
  assign b_i_k_0_i_j_8 = _T_2462;	// matmul/matmul-hw.mlir:18866:5
  //PROBE: b_i_k_0_i_j_8	// matmul/matmul-hw.mlir:18867:5
  assign c_prev_i_k_0_i_j_8 = C_reg_bank0_p0_rd_data_2317;	// matmul/matmul-hw.mlir:18839:36, :18869:5
  //PROBE: c_prev_i_k_0_i_j_8	// matmul/matmul-hw.mlir:18870:5
  assign tk_i_k_0_i_j_8 = _T_2797;	// matmul/matmul-hw.mlir:18872:5
  //PROBE: tk_i_k_0_i_j_8	// matmul/matmul-hw.mlir:18873:5
  wire [31:0] _T_3497 = mult_inst128_result + C_reg_bank0_p0_rd_data_2317;	// matmul/matmul-hw.mlir:18839:36, :18860:28, :18874:13
  assign c_i_k_0_i_j_8 = _T_3497;	// matmul/matmul-hw.mlir:18876:5
  //PROBE: c_i_k_0_i_j_8	// matmul/matmul-hw.mlir:18877:5
  assign _T_689 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18878:13
  assign _T_688 = _T_2841 ? _T_3497 : 32'bx;	// matmul/matmul-hw.mlir:8723:19, :18879:13
  localparam [3:0] _T_3499 = 4'h0;	// matmul/matmul-hw.mlir:18882:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18883:5
    if (rst)	// matmul/matmul-hw.mlir:18883:5
      i_k_next_3498 <= _T_3499;	// matmul/matmul-hw.mlir:18886:7
    else	// matmul/matmul-hw.mlir:18883:5
      i_k_next_3498 <= i_j_next_3478;	// matmul/matmul-hw.mlir:18764:13, :18884:7
  end // always @(posedge)
  assign _T_687 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18888:13
  assign _T_686 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18889:13
  mult mult_inst129 (	// matmul/matmul-hw.mlir:18890:28
    .a      (A_reg_bank129_p0_rd_data),	// matmul/matmul-hw.mlir:12344:33
    .b      (_T_2478),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst129_result)
  );
  assign _T_685 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18891:13
  assign a_i_k_1_i_j_8 = A_reg_bank129_p0_rd_data;	// matmul/matmul-hw.mlir:12344:33, :18893:5
  //PROBE: a_i_k_1_i_j_8	// matmul/matmul-hw.mlir:18894:5
  assign b_i_k_1_i_j_8 = _T_2478;	// matmul/matmul-hw.mlir:18896:5
  //PROBE: b_i_k_1_i_j_8	// matmul/matmul-hw.mlir:18897:5
  assign c_prev_i_k_1_i_j_8 = C_reg_bank1_p0_rd_data_2316;	// matmul/matmul-hw.mlir:18840:36, :18899:5
  //PROBE: c_prev_i_k_1_i_j_8	// matmul/matmul-hw.mlir:18900:5
  assign tk_i_k_1_i_j_8 = _T_2808;	// matmul/matmul-hw.mlir:18902:5
  //PROBE: tk_i_k_1_i_j_8	// matmul/matmul-hw.mlir:18903:5
  wire [31:0] _T_3500 = mult_inst129_result + C_reg_bank1_p0_rd_data_2316;	// matmul/matmul-hw.mlir:18840:36, :18890:28, :18904:13
  assign c_i_k_1_i_j_8 = _T_3500;	// matmul/matmul-hw.mlir:18906:5
  //PROBE: c_i_k_1_i_j_8	// matmul/matmul-hw.mlir:18907:5
  assign _T_684 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18908:13
  assign _T_683 = _T_2852 ? _T_3500 : 32'bx;	// matmul/matmul-hw.mlir:8718:19, :18909:13
  localparam [3:0] _T_3502 = 4'h0;	// matmul/matmul-hw.mlir:18912:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18913:5
    if (rst)	// matmul/matmul-hw.mlir:18913:5
      i_k_next_3501 <= _T_3502;	// matmul/matmul-hw.mlir:18916:7
    else	// matmul/matmul-hw.mlir:18913:5
      i_k_next_3501 <= i_k_next_3498;	// matmul/matmul-hw.mlir:18881:13, :18914:7
  end // always @(posedge)
  assign _T_682 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18918:13
  assign _T_681 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18919:13
  mult mult_inst130 (	// matmul/matmul-hw.mlir:18920:28
    .a      (A_reg_bank130_p0_rd_data),	// matmul/matmul-hw.mlir:12345:33
    .b      (_T_2494),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst130_result)
  );
  assign _T_680 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18921:13
  assign a_i_k_2_i_j_8 = A_reg_bank130_p0_rd_data;	// matmul/matmul-hw.mlir:12345:33, :18923:5
  //PROBE: a_i_k_2_i_j_8	// matmul/matmul-hw.mlir:18924:5
  assign b_i_k_2_i_j_8 = _T_2494;	// matmul/matmul-hw.mlir:18926:5
  //PROBE: b_i_k_2_i_j_8	// matmul/matmul-hw.mlir:18927:5
  assign c_prev_i_k_2_i_j_8 = C_reg_bank2_p0_rd_data_2315;	// matmul/matmul-hw.mlir:18841:36, :18929:5
  //PROBE: c_prev_i_k_2_i_j_8	// matmul/matmul-hw.mlir:18930:5
  assign tk_i_k_2_i_j_8 = _T_2819;	// matmul/matmul-hw.mlir:18932:5
  //PROBE: tk_i_k_2_i_j_8	// matmul/matmul-hw.mlir:18933:5
  wire [31:0] _T_3503 = mult_inst130_result + C_reg_bank2_p0_rd_data_2315;	// matmul/matmul-hw.mlir:18841:36, :18920:28, :18934:13
  assign c_i_k_2_i_j_8 = _T_3503;	// matmul/matmul-hw.mlir:18936:5
  //PROBE: c_i_k_2_i_j_8	// matmul/matmul-hw.mlir:18937:5
  assign _T_679 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18938:13
  assign _T_678 = _T_2863 ? _T_3503 : 32'bx;	// matmul/matmul-hw.mlir:8713:19, :18939:13
  localparam [3:0] _T_3505 = 4'h0;	// matmul/matmul-hw.mlir:18942:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18943:5
    if (rst)	// matmul/matmul-hw.mlir:18943:5
      i_k_next_3504 <= _T_3505;	// matmul/matmul-hw.mlir:18946:7
    else	// matmul/matmul-hw.mlir:18943:5
      i_k_next_3504 <= i_k_next_3501;	// matmul/matmul-hw.mlir:18911:13, :18944:7
  end // always @(posedge)
  assign _T_677 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18948:13
  assign _T_676 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18949:13
  mult mult_inst131 (	// matmul/matmul-hw.mlir:18950:28
    .a      (A_reg_bank131_p0_rd_data),	// matmul/matmul-hw.mlir:12346:33
    .b      (_T_2510),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst131_result)
  );
  assign _T_675 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18951:13
  assign a_i_k_3_i_j_8 = A_reg_bank131_p0_rd_data;	// matmul/matmul-hw.mlir:12346:33, :18953:5
  //PROBE: a_i_k_3_i_j_8	// matmul/matmul-hw.mlir:18954:5
  assign b_i_k_3_i_j_8 = _T_2510;	// matmul/matmul-hw.mlir:18956:5
  //PROBE: b_i_k_3_i_j_8	// matmul/matmul-hw.mlir:18957:5
  assign c_prev_i_k_3_i_j_8 = C_reg_bank3_p0_rd_data_2314;	// matmul/matmul-hw.mlir:18842:36, :18959:5
  //PROBE: c_prev_i_k_3_i_j_8	// matmul/matmul-hw.mlir:18960:5
  assign tk_i_k_3_i_j_8 = _T_2830;	// matmul/matmul-hw.mlir:18962:5
  //PROBE: tk_i_k_3_i_j_8	// matmul/matmul-hw.mlir:18963:5
  wire [31:0] _T_3506 = mult_inst131_result + C_reg_bank3_p0_rd_data_2314;	// matmul/matmul-hw.mlir:18842:36, :18950:28, :18964:13
  assign c_i_k_3_i_j_8 = _T_3506;	// matmul/matmul-hw.mlir:18966:5
  //PROBE: c_i_k_3_i_j_8	// matmul/matmul-hw.mlir:18967:5
  assign _T_674 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18968:13
  assign _T_673 = _T_2874 ? _T_3506 : 32'bx;	// matmul/matmul-hw.mlir:8708:19, :18969:13
  localparam [3:0] _T_3508 = 4'h0;	// matmul/matmul-hw.mlir:18972:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:18973:5
    if (rst)	// matmul/matmul-hw.mlir:18973:5
      i_k_next_3507 <= _T_3508;	// matmul/matmul-hw.mlir:18976:7
    else	// matmul/matmul-hw.mlir:18973:5
      i_k_next_3507 <= i_k_next_3504;	// matmul/matmul-hw.mlir:18941:13, :18974:7
  end // always @(posedge)
  assign _T_672 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18978:13
  assign _T_671 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18979:13
  mult mult_inst132 (	// matmul/matmul-hw.mlir:18980:28
    .a      (A_reg_bank132_p0_rd_data),	// matmul/matmul-hw.mlir:12347:33
    .b      (_T_2526),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst132_result)
  );
  assign _T_670 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18981:13
  assign a_i_k_4_i_j_8 = A_reg_bank132_p0_rd_data;	// matmul/matmul-hw.mlir:12347:33, :18983:5
  //PROBE: a_i_k_4_i_j_8	// matmul/matmul-hw.mlir:18984:5
  assign b_i_k_4_i_j_8 = _T_2526;	// matmul/matmul-hw.mlir:18986:5
  //PROBE: b_i_k_4_i_j_8	// matmul/matmul-hw.mlir:18987:5
  assign c_prev_i_k_4_i_j_8 = C_reg_bank4_p0_rd_data_2313;	// matmul/matmul-hw.mlir:18843:36, :18989:5
  //PROBE: c_prev_i_k_4_i_j_8	// matmul/matmul-hw.mlir:18990:5
  assign tk_i_k_4_i_j_8 = _T_2841;	// matmul/matmul-hw.mlir:18992:5
  //PROBE: tk_i_k_4_i_j_8	// matmul/matmul-hw.mlir:18993:5
  wire [31:0] _T_3509 = mult_inst132_result + C_reg_bank4_p0_rd_data_2313;	// matmul/matmul-hw.mlir:18843:36, :18980:28, :18994:13
  assign c_i_k_4_i_j_8 = _T_3509;	// matmul/matmul-hw.mlir:18996:5
  //PROBE: c_i_k_4_i_j_8	// matmul/matmul-hw.mlir:18997:5
  assign _T_669 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :18998:13
  assign _T_668 = _T_2885 ? _T_3509 : 32'bx;	// matmul/matmul-hw.mlir:8703:19, :18999:13
  localparam [3:0] _T_3511 = 4'h0;	// matmul/matmul-hw.mlir:19002:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19003:5
    if (rst)	// matmul/matmul-hw.mlir:19003:5
      i_k_next_3510 <= _T_3511;	// matmul/matmul-hw.mlir:19006:7
    else	// matmul/matmul-hw.mlir:19003:5
      i_k_next_3510 <= i_k_next_3507;	// matmul/matmul-hw.mlir:18971:13, :19004:7
  end // always @(posedge)
  assign _T_667 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19008:13
  assign _T_666 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19009:13
  mult mult_inst133 (	// matmul/matmul-hw.mlir:19010:28
    .a      (A_reg_bank133_p0_rd_data),	// matmul/matmul-hw.mlir:12348:33
    .b      (_T_2542),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst133_result)
  );
  assign _T_665 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19011:13
  assign a_i_k_5_i_j_8 = A_reg_bank133_p0_rd_data;	// matmul/matmul-hw.mlir:12348:33, :19013:5
  //PROBE: a_i_k_5_i_j_8	// matmul/matmul-hw.mlir:19014:5
  assign b_i_k_5_i_j_8 = _T_2542;	// matmul/matmul-hw.mlir:19016:5
  //PROBE: b_i_k_5_i_j_8	// matmul/matmul-hw.mlir:19017:5
  assign c_prev_i_k_5_i_j_8 = C_reg_bank5_p0_rd_data_2312;	// matmul/matmul-hw.mlir:18844:36, :19019:5
  //PROBE: c_prev_i_k_5_i_j_8	// matmul/matmul-hw.mlir:19020:5
  assign tk_i_k_5_i_j_8 = _T_2852;	// matmul/matmul-hw.mlir:19022:5
  //PROBE: tk_i_k_5_i_j_8	// matmul/matmul-hw.mlir:19023:5
  wire [31:0] _T_3512 = mult_inst133_result + C_reg_bank5_p0_rd_data_2312;	// matmul/matmul-hw.mlir:18844:36, :19010:28, :19024:13
  assign c_i_k_5_i_j_8 = _T_3512;	// matmul/matmul-hw.mlir:19026:5
  //PROBE: c_i_k_5_i_j_8	// matmul/matmul-hw.mlir:19027:5
  assign _T_664 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19028:13
  assign _T_663 = _T_2892 ? _T_3512 : 32'bx;	// matmul/matmul-hw.mlir:8698:19, :19029:13
  localparam [3:0] _T_3514 = 4'h0;	// matmul/matmul-hw.mlir:19032:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19033:5
    if (rst)	// matmul/matmul-hw.mlir:19033:5
      i_k_next_3513 <= _T_3514;	// matmul/matmul-hw.mlir:19036:7
    else	// matmul/matmul-hw.mlir:19033:5
      i_k_next_3513 <= i_k_next_3510;	// matmul/matmul-hw.mlir:19001:13, :19034:7
  end // always @(posedge)
  assign _T_662 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19038:13
  assign _T_661 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19039:13
  mult mult_inst134 (	// matmul/matmul-hw.mlir:19040:28
    .a      (A_reg_bank134_p0_rd_data),	// matmul/matmul-hw.mlir:12349:33
    .b      (_T_2558),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst134_result)
  );
  assign _T_660 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19041:13
  assign a_i_k_6_i_j_8 = A_reg_bank134_p0_rd_data;	// matmul/matmul-hw.mlir:12349:33, :19043:5
  //PROBE: a_i_k_6_i_j_8	// matmul/matmul-hw.mlir:19044:5
  assign b_i_k_6_i_j_8 = _T_2558;	// matmul/matmul-hw.mlir:19046:5
  //PROBE: b_i_k_6_i_j_8	// matmul/matmul-hw.mlir:19047:5
  assign c_prev_i_k_6_i_j_8 = C_reg_bank6_p0_rd_data_2311;	// matmul/matmul-hw.mlir:18845:36, :19049:5
  //PROBE: c_prev_i_k_6_i_j_8	// matmul/matmul-hw.mlir:19050:5
  assign tk_i_k_6_i_j_8 = _T_2863;	// matmul/matmul-hw.mlir:19052:5
  //PROBE: tk_i_k_6_i_j_8	// matmul/matmul-hw.mlir:19053:5
  wire [31:0] _T_3515 = mult_inst134_result + C_reg_bank6_p0_rd_data_2311;	// matmul/matmul-hw.mlir:18845:36, :19040:28, :19054:13
  assign c_i_k_6_i_j_8 = _T_3515;	// matmul/matmul-hw.mlir:19056:5
  //PROBE: c_i_k_6_i_j_8	// matmul/matmul-hw.mlir:19057:5
  assign _T_659 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19058:13
  assign _T_658 = _T_2897 ? _T_3515 : 32'bx;	// matmul/matmul-hw.mlir:8693:19, :19059:13
  localparam [3:0] _T_3517 = 4'h0;	// matmul/matmul-hw.mlir:19062:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19063:5
    if (rst)	// matmul/matmul-hw.mlir:19063:5
      i_k_next_3516 <= _T_3517;	// matmul/matmul-hw.mlir:19066:7
    else	// matmul/matmul-hw.mlir:19063:5
      i_k_next_3516 <= i_k_next_3513;	// matmul/matmul-hw.mlir:19031:13, :19064:7
  end // always @(posedge)
  assign _T_657 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19068:13
  assign _T_656 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19069:13
  mult mult_inst135 (	// matmul/matmul-hw.mlir:19070:28
    .a      (A_reg_bank135_p0_rd_data),	// matmul/matmul-hw.mlir:12350:33
    .b      (_T_2574),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst135_result)
  );
  assign _T_655 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19071:13
  assign a_i_k_7_i_j_8 = A_reg_bank135_p0_rd_data;	// matmul/matmul-hw.mlir:12350:33, :19073:5
  //PROBE: a_i_k_7_i_j_8	// matmul/matmul-hw.mlir:19074:5
  assign b_i_k_7_i_j_8 = _T_2574;	// matmul/matmul-hw.mlir:19076:5
  //PROBE: b_i_k_7_i_j_8	// matmul/matmul-hw.mlir:19077:5
  assign c_prev_i_k_7_i_j_8 = C_reg_bank7_p0_rd_data_2310;	// matmul/matmul-hw.mlir:18846:36, :19079:5
  //PROBE: c_prev_i_k_7_i_j_8	// matmul/matmul-hw.mlir:19080:5
  assign tk_i_k_7_i_j_8 = _T_2874;	// matmul/matmul-hw.mlir:19082:5
  //PROBE: tk_i_k_7_i_j_8	// matmul/matmul-hw.mlir:19083:5
  wire [31:0] _T_3518 = mult_inst135_result + C_reg_bank7_p0_rd_data_2310;	// matmul/matmul-hw.mlir:18846:36, :19070:28, :19084:13
  assign c_i_k_7_i_j_8 = _T_3518;	// matmul/matmul-hw.mlir:19086:5
  //PROBE: c_i_k_7_i_j_8	// matmul/matmul-hw.mlir:19087:5
  assign _T_654 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19088:13
  assign _T_653 = _T_2902 ? _T_3518 : 32'bx;	// matmul/matmul-hw.mlir:8688:19, :19089:13
  localparam [3:0] _T_3520 = 4'h0;	// matmul/matmul-hw.mlir:19092:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19093:5
    if (rst)	// matmul/matmul-hw.mlir:19093:5
      i_k_next_3519 <= _T_3520;	// matmul/matmul-hw.mlir:19096:7
    else	// matmul/matmul-hw.mlir:19093:5
      i_k_next_3519 <= i_k_next_3516;	// matmul/matmul-hw.mlir:19061:13, :19094:7
  end // always @(posedge)
  assign _T_652 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19098:13
  assign _T_651 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19099:13
  mult mult_inst136 (	// matmul/matmul-hw.mlir:19100:28
    .a      (A_reg_bank136_p0_rd_data),	// matmul/matmul-hw.mlir:12351:33
    .b      (_T_2590),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst136_result)
  );
  assign _T_650 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19101:13
  assign a_i_k_8_i_j_8 = A_reg_bank136_p0_rd_data;	// matmul/matmul-hw.mlir:12351:33, :19103:5
  //PROBE: a_i_k_8_i_j_8	// matmul/matmul-hw.mlir:19104:5
  assign b_i_k_8_i_j_8 = _T_2590;	// matmul/matmul-hw.mlir:19106:5
  //PROBE: b_i_k_8_i_j_8	// matmul/matmul-hw.mlir:19107:5
  assign c_prev_i_k_8_i_j_8 = C_reg_bank8_p0_rd_data_2309;	// matmul/matmul-hw.mlir:18847:36, :19109:5
  //PROBE: c_prev_i_k_8_i_j_8	// matmul/matmul-hw.mlir:19110:5
  assign tk_i_k_8_i_j_8 = _T_2885;	// matmul/matmul-hw.mlir:19112:5
  //PROBE: tk_i_k_8_i_j_8	// matmul/matmul-hw.mlir:19113:5
  wire [31:0] _T_3521 = mult_inst136_result + C_reg_bank8_p0_rd_data_2309;	// matmul/matmul-hw.mlir:18847:36, :19100:28, :19114:13
  assign c_i_k_8_i_j_8 = _T_3521;	// matmul/matmul-hw.mlir:19116:5
  //PROBE: c_i_k_8_i_j_8	// matmul/matmul-hw.mlir:19117:5
  assign _T_649 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19118:13
  assign _T_648 = _T_2907 ? _T_3521 : 32'bx;	// matmul/matmul-hw.mlir:8683:19, :19119:13
  localparam [3:0] _T_3523 = 4'h0;	// matmul/matmul-hw.mlir:19122:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19123:5
    if (rst)	// matmul/matmul-hw.mlir:19123:5
      i_k_next_3522 <= _T_3523;	// matmul/matmul-hw.mlir:19126:7
    else	// matmul/matmul-hw.mlir:19123:5
      i_k_next_3522 <= i_k_next_3519;	// matmul/matmul-hw.mlir:19091:13, :19124:7
  end // always @(posedge)
  assign _T_647 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19128:13
  assign _T_646 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19129:13
  mult mult_inst137 (	// matmul/matmul-hw.mlir:19130:28
    .a      (A_reg_bank137_p0_rd_data),	// matmul/matmul-hw.mlir:12352:33
    .b      (_T_2606),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst137_result)
  );
  assign _T_645 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19131:13
  assign a_i_k_9_i_j_8 = A_reg_bank137_p0_rd_data;	// matmul/matmul-hw.mlir:12352:33, :19133:5
  //PROBE: a_i_k_9_i_j_8	// matmul/matmul-hw.mlir:19134:5
  assign b_i_k_9_i_j_8 = _T_2606;	// matmul/matmul-hw.mlir:19136:5
  //PROBE: b_i_k_9_i_j_8	// matmul/matmul-hw.mlir:19137:5
  assign c_prev_i_k_9_i_j_8 = C_reg_bank9_p0_rd_data_2308;	// matmul/matmul-hw.mlir:18848:36, :19139:5
  //PROBE: c_prev_i_k_9_i_j_8	// matmul/matmul-hw.mlir:19140:5
  assign tk_i_k_9_i_j_8 = _T_2892;	// matmul/matmul-hw.mlir:19142:5
  //PROBE: tk_i_k_9_i_j_8	// matmul/matmul-hw.mlir:19143:5
  wire [31:0] _T_3524 = mult_inst137_result + C_reg_bank9_p0_rd_data_2308;	// matmul/matmul-hw.mlir:18848:36, :19130:28, :19144:13
  assign c_i_k_9_i_j_8 = _T_3524;	// matmul/matmul-hw.mlir:19146:5
  //PROBE: c_i_k_9_i_j_8	// matmul/matmul-hw.mlir:19147:5
  assign _T_644 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19148:13
  assign _T_643 = _T_2912 ? _T_3524 : 32'bx;	// matmul/matmul-hw.mlir:8678:19, :19149:13
  localparam [3:0] _T_3526 = 4'h0;	// matmul/matmul-hw.mlir:19152:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19153:5
    if (rst)	// matmul/matmul-hw.mlir:19153:5
      i_k_next_3525 <= _T_3526;	// matmul/matmul-hw.mlir:19156:7
    else	// matmul/matmul-hw.mlir:19153:5
      i_k_next_3525 <= i_k_next_3522;	// matmul/matmul-hw.mlir:19121:13, :19154:7
  end // always @(posedge)
  assign _T_642 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19158:13
  assign _T_641 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19159:13
  mult mult_inst138 (	// matmul/matmul-hw.mlir:19160:28
    .a      (A_reg_bank138_p0_rd_data),	// matmul/matmul-hw.mlir:12353:33
    .b      (_T_2622),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst138_result)
  );
  assign _T_640 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19161:13
  assign a_i_k_10_i_j_8 = A_reg_bank138_p0_rd_data;	// matmul/matmul-hw.mlir:12353:33, :19163:5
  //PROBE: a_i_k_10_i_j_8	// matmul/matmul-hw.mlir:19164:5
  assign b_i_k_10_i_j_8 = _T_2622;	// matmul/matmul-hw.mlir:19166:5
  //PROBE: b_i_k_10_i_j_8	// matmul/matmul-hw.mlir:19167:5
  assign c_prev_i_k_10_i_j_8 = C_reg_bank10_p0_rd_data_2307;	// matmul/matmul-hw.mlir:18849:37, :19169:5
  //PROBE: c_prev_i_k_10_i_j_8	// matmul/matmul-hw.mlir:19170:5
  assign tk_i_k_10_i_j_8 = _T_2897;	// matmul/matmul-hw.mlir:19172:5
  //PROBE: tk_i_k_10_i_j_8	// matmul/matmul-hw.mlir:19173:5
  wire [31:0] _T_3527 = mult_inst138_result + C_reg_bank10_p0_rd_data_2307;	// matmul/matmul-hw.mlir:18849:37, :19160:28, :19174:13
  assign c_i_k_10_i_j_8 = _T_3527;	// matmul/matmul-hw.mlir:19176:5
  //PROBE: c_i_k_10_i_j_8	// matmul/matmul-hw.mlir:19177:5
  assign _T_639 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19178:13
  assign _T_638 = _T_2917 ? _T_3527 : 32'bx;	// matmul/matmul-hw.mlir:8673:19, :19179:13
  localparam [3:0] _T_3529 = 4'h0;	// matmul/matmul-hw.mlir:19182:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19183:5
    if (rst)	// matmul/matmul-hw.mlir:19183:5
      i_k_next_3528 <= _T_3529;	// matmul/matmul-hw.mlir:19186:7
    else	// matmul/matmul-hw.mlir:19183:5
      i_k_next_3528 <= i_k_next_3525;	// matmul/matmul-hw.mlir:19151:13, :19184:7
  end // always @(posedge)
  assign _T_637 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19188:13
  assign _T_636 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19189:13
  mult mult_inst139 (	// matmul/matmul-hw.mlir:19190:28
    .a      (A_reg_bank139_p0_rd_data),	// matmul/matmul-hw.mlir:12354:33
    .b      (_T_2638),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst139_result)
  );
  assign _T_635 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19191:13
  assign a_i_k_11_i_j_8 = A_reg_bank139_p0_rd_data;	// matmul/matmul-hw.mlir:12354:33, :19193:5
  //PROBE: a_i_k_11_i_j_8	// matmul/matmul-hw.mlir:19194:5
  assign b_i_k_11_i_j_8 = _T_2638;	// matmul/matmul-hw.mlir:19196:5
  //PROBE: b_i_k_11_i_j_8	// matmul/matmul-hw.mlir:19197:5
  assign c_prev_i_k_11_i_j_8 = C_reg_bank11_p0_rd_data_2306;	// matmul/matmul-hw.mlir:18850:37, :19199:5
  //PROBE: c_prev_i_k_11_i_j_8	// matmul/matmul-hw.mlir:19200:5
  assign tk_i_k_11_i_j_8 = _T_2902;	// matmul/matmul-hw.mlir:19202:5
  //PROBE: tk_i_k_11_i_j_8	// matmul/matmul-hw.mlir:19203:5
  wire [31:0] _T_3530 = mult_inst139_result + C_reg_bank11_p0_rd_data_2306;	// matmul/matmul-hw.mlir:18850:37, :19190:28, :19204:13
  assign c_i_k_11_i_j_8 = _T_3530;	// matmul/matmul-hw.mlir:19206:5
  //PROBE: c_i_k_11_i_j_8	// matmul/matmul-hw.mlir:19207:5
  assign _T_634 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19208:13
  assign _T_633 = _T_2922 ? _T_3530 : 32'bx;	// matmul/matmul-hw.mlir:8668:18, :19209:13
  localparam [3:0] _T_3532 = 4'h0;	// matmul/matmul-hw.mlir:19212:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19213:5
    if (rst)	// matmul/matmul-hw.mlir:19213:5
      i_k_next_3531 <= _T_3532;	// matmul/matmul-hw.mlir:19216:7
    else	// matmul/matmul-hw.mlir:19213:5
      i_k_next_3531 <= i_k_next_3528;	// matmul/matmul-hw.mlir:19181:13, :19214:7
  end // always @(posedge)
  assign _T_632 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19218:13
  assign _T_631 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19219:13
  mult mult_inst140 (	// matmul/matmul-hw.mlir:19220:28
    .a      (A_reg_bank140_p0_rd_data),	// matmul/matmul-hw.mlir:12355:33
    .b      (_T_2654),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst140_result)
  );
  assign _T_630 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19221:13
  assign a_i_k_12_i_j_8 = A_reg_bank140_p0_rd_data;	// matmul/matmul-hw.mlir:12355:33, :19223:5
  //PROBE: a_i_k_12_i_j_8	// matmul/matmul-hw.mlir:19224:5
  assign b_i_k_12_i_j_8 = _T_2654;	// matmul/matmul-hw.mlir:19226:5
  //PROBE: b_i_k_12_i_j_8	// matmul/matmul-hw.mlir:19227:5
  assign c_prev_i_k_12_i_j_8 = C_reg_bank12_p0_rd_data_2305;	// matmul/matmul-hw.mlir:18851:37, :19229:5
  //PROBE: c_prev_i_k_12_i_j_8	// matmul/matmul-hw.mlir:19230:5
  assign tk_i_k_12_i_j_8 = _T_2907;	// matmul/matmul-hw.mlir:19232:5
  //PROBE: tk_i_k_12_i_j_8	// matmul/matmul-hw.mlir:19233:5
  wire [31:0] _T_3533 = mult_inst140_result + C_reg_bank12_p0_rd_data_2305;	// matmul/matmul-hw.mlir:18851:37, :19220:28, :19234:13
  assign c_i_k_12_i_j_8 = _T_3533;	// matmul/matmul-hw.mlir:19236:5
  //PROBE: c_i_k_12_i_j_8	// matmul/matmul-hw.mlir:19237:5
  assign _T_629 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19238:13
  assign _T_628 = _T_2927 ? _T_3533 : 32'bx;	// matmul/matmul-hw.mlir:8663:18, :19239:13
  localparam [3:0] _T_3535 = 4'h0;	// matmul/matmul-hw.mlir:19242:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19243:5
    if (rst)	// matmul/matmul-hw.mlir:19243:5
      i_k_next_3534 <= _T_3535;	// matmul/matmul-hw.mlir:19246:7
    else	// matmul/matmul-hw.mlir:19243:5
      i_k_next_3534 <= i_k_next_3531;	// matmul/matmul-hw.mlir:19211:13, :19244:7
  end // always @(posedge)
  assign _T_627 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19248:13
  assign _T_626 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19249:13
  mult mult_inst141 (	// matmul/matmul-hw.mlir:19250:28
    .a      (A_reg_bank141_p0_rd_data),	// matmul/matmul-hw.mlir:12356:33
    .b      (_T_2670),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst141_result)
  );
  assign _T_625 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19251:13
  assign a_i_k_13_i_j_8 = A_reg_bank141_p0_rd_data;	// matmul/matmul-hw.mlir:12356:33, :19253:5
  //PROBE: a_i_k_13_i_j_8	// matmul/matmul-hw.mlir:19254:5
  assign b_i_k_13_i_j_8 = _T_2670;	// matmul/matmul-hw.mlir:19256:5
  //PROBE: b_i_k_13_i_j_8	// matmul/matmul-hw.mlir:19257:5
  assign c_prev_i_k_13_i_j_8 = C_reg_bank13_p0_rd_data_2304;	// matmul/matmul-hw.mlir:18852:37, :19259:5
  //PROBE: c_prev_i_k_13_i_j_8	// matmul/matmul-hw.mlir:19260:5
  assign tk_i_k_13_i_j_8 = _T_2912;	// matmul/matmul-hw.mlir:19262:5
  //PROBE: tk_i_k_13_i_j_8	// matmul/matmul-hw.mlir:19263:5
  wire [31:0] _T_3536 = mult_inst141_result + C_reg_bank13_p0_rd_data_2304;	// matmul/matmul-hw.mlir:18852:37, :19250:28, :19264:13
  assign c_i_k_13_i_j_8 = _T_3536;	// matmul/matmul-hw.mlir:19266:5
  //PROBE: c_i_k_13_i_j_8	// matmul/matmul-hw.mlir:19267:5
  assign _T_624 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19268:13
  assign _T_623 = _T_2932 ? _T_3536 : 32'bx;	// matmul/matmul-hw.mlir:8658:18, :19269:13
  localparam [3:0] _T_3538 = 4'h0;	// matmul/matmul-hw.mlir:19272:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19273:5
    if (rst)	// matmul/matmul-hw.mlir:19273:5
      i_k_next_3537 <= _T_3538;	// matmul/matmul-hw.mlir:19276:7
    else	// matmul/matmul-hw.mlir:19273:5
      i_k_next_3537 <= i_k_next_3534;	// matmul/matmul-hw.mlir:19241:13, :19274:7
  end // always @(posedge)
  assign _T_622 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19278:13
  assign _T_621 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19279:13
  mult mult_inst142 (	// matmul/matmul-hw.mlir:19280:28
    .a      (A_reg_bank142_p0_rd_data),	// matmul/matmul-hw.mlir:12357:33
    .b      (_T_2686),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst142_result)
  );
  assign _T_620 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19281:13
  assign a_i_k_14_i_j_8 = A_reg_bank142_p0_rd_data;	// matmul/matmul-hw.mlir:12357:33, :19283:5
  //PROBE: a_i_k_14_i_j_8	// matmul/matmul-hw.mlir:19284:5
  assign b_i_k_14_i_j_8 = _T_2686;	// matmul/matmul-hw.mlir:19286:5
  //PROBE: b_i_k_14_i_j_8	// matmul/matmul-hw.mlir:19287:5
  assign c_prev_i_k_14_i_j_8 = C_reg_bank14_p0_rd_data_2303;	// matmul/matmul-hw.mlir:18853:37, :19289:5
  //PROBE: c_prev_i_k_14_i_j_8	// matmul/matmul-hw.mlir:19290:5
  assign tk_i_k_14_i_j_8 = _T_2917;	// matmul/matmul-hw.mlir:19292:5
  //PROBE: tk_i_k_14_i_j_8	// matmul/matmul-hw.mlir:19293:5
  wire [31:0] _T_3539 = mult_inst142_result + C_reg_bank14_p0_rd_data_2303;	// matmul/matmul-hw.mlir:18853:37, :19280:28, :19294:13
  assign c_i_k_14_i_j_8 = _T_3539;	// matmul/matmul-hw.mlir:19296:5
  //PROBE: c_i_k_14_i_j_8	// matmul/matmul-hw.mlir:19297:5
  assign _T_619 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19298:13
  assign _T_618 = _T_2937 ? _T_3539 : 32'bx;	// matmul/matmul-hw.mlir:8653:18, :19299:13
  localparam [3:0] _T_3541 = 4'h0;	// matmul/matmul-hw.mlir:19302:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19303:5
    if (rst)	// matmul/matmul-hw.mlir:19303:5
      i_k_next_3540 <= _T_3541;	// matmul/matmul-hw.mlir:19306:7
    else	// matmul/matmul-hw.mlir:19303:5
      i_k_next_3540 <= i_k_next_3537;	// matmul/matmul-hw.mlir:19271:13, :19304:7
  end // always @(posedge)
  assign _T_617 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19308:13
  assign _T_616 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19309:13
  mult mult_inst143 (	// matmul/matmul-hw.mlir:19310:28
    .a      (A_reg_bank143_p0_rd_data),	// matmul/matmul-hw.mlir:12358:33
    .b      (_T_2702),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst143_result)
  );
  assign _T_615 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19311:13
  assign a_i_k_15_i_j_8 = A_reg_bank143_p0_rd_data;	// matmul/matmul-hw.mlir:12358:33, :19313:5
  //PROBE: a_i_k_15_i_j_8	// matmul/matmul-hw.mlir:19314:5
  assign b_i_k_15_i_j_8 = _T_2702;	// matmul/matmul-hw.mlir:19316:5
  //PROBE: b_i_k_15_i_j_8	// matmul/matmul-hw.mlir:19317:5
  assign c_prev_i_k_15_i_j_8 = C_reg_bank15_p0_rd_data_2302;	// matmul/matmul-hw.mlir:18854:37, :19319:5
  //PROBE: c_prev_i_k_15_i_j_8	// matmul/matmul-hw.mlir:19320:5
  assign tk_i_k_15_i_j_8 = _T_2922;	// matmul/matmul-hw.mlir:19322:5
  //PROBE: tk_i_k_15_i_j_8	// matmul/matmul-hw.mlir:19323:5
  wire [31:0] _T_3542 = mult_inst143_result + C_reg_bank15_p0_rd_data_2302;	// matmul/matmul-hw.mlir:18854:37, :19310:28, :19324:13
  assign c_i_k_15_i_j_8 = _T_3542;	// matmul/matmul-hw.mlir:19326:5
  //PROBE: c_i_k_15_i_j_8	// matmul/matmul-hw.mlir:19327:5
  assign _T_614 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19328:13
  assign _T_613 = _T_2942 ? _T_3542 : 32'bx;	// matmul/matmul-hw.mlir:8648:18, :19329:13
  localparam [3:0] _T_3544 = 4'h0;	// matmul/matmul-hw.mlir:19332:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19333:5
    if (rst)	// matmul/matmul-hw.mlir:19333:5
      i_k_next_3543 <= _T_3544;	// matmul/matmul-hw.mlir:19336:7
    else	// matmul/matmul-hw.mlir:19333:5
      i_k_next_3543 <= i_k_next_3540;	// matmul/matmul-hw.mlir:19301:13, :19334:7
  end // always @(posedge)
  assign _T_612 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19338:13
  wire [3:0][3:0] _T_3546 = i_delayed_3545;	// matmul/matmul-hw.mlir:19340:13
  wire [3:0][3:0] _T_3547 = {_T_3546[2'h0+:3], {{i_k_next_3543}}};	// matmul/matmul-hw.mlir:19331:13, :19341:19, :19342:13, :19343:13, :19344:13
  wire [3:0][3:0] _T_3548 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:19345:19, :19346:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19347:5
    if (rst)	// matmul/matmul-hw.mlir:19347:5
      i_delayed_3545 <= _T_3548;	// matmul/matmul-hw.mlir:19350:7
    else	// matmul/matmul-hw.mlir:19347:5
      i_delayed_3545 <= _T_3547;	// matmul/matmul-hw.mlir:19348:7
  end // always @(posedge)
  assign _T_611 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19354:13
  assign _T_610 = _T_2947 ? i_delayed_3545[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8645:17, :19340:13, :19352:20, :19353:13, :19355:13
  assign _T_609 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19356:13
  assign _T_608 = _T_2947 ? C_reg_bank16_p0_rd_data_2301 : 32'bx;	// matmul/matmul-hw.mlir:8643:18, :18855:37, :19357:13
  localparam [3:0] _T_3550 = 4'h0;	// matmul/matmul-hw.mlir:19360:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19361:5
    if (rst)	// matmul/matmul-hw.mlir:19361:5
      i_j_next_3549 <= _T_3550;	// matmul/matmul-hw.mlir:19364:7
    else	// matmul/matmul-hw.mlir:19361:5
      i_j_next_3549 <= i_j_next_3478;	// matmul/matmul-hw.mlir:18764:13, :19362:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3551 (	// matmul/matmul-hw.mlir:19434:36
    .p0_rd_en   (_T_603),	// matmul/matmul-hw.mlir:19456:13
    .p1_wr_en   (_T_607),	// matmul/matmul-hw.mlir:19451:13
    .p1_wr_data (_T_606),	// matmul/matmul-hw.mlir:19452:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2300)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3552 (	// matmul/matmul-hw.mlir:19435:36
    .p0_rd_en   (_T_598),	// matmul/matmul-hw.mlir:19486:13
    .p1_wr_en   (_T_602),	// matmul/matmul-hw.mlir:19473:13
    .p1_wr_data (_T_601),	// matmul/matmul-hw.mlir:19474:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2299)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3553 (	// matmul/matmul-hw.mlir:19436:36
    .p0_rd_en   (_T_593),	// matmul/matmul-hw.mlir:19516:13
    .p1_wr_en   (_T_597),	// matmul/matmul-hw.mlir:19503:13
    .p1_wr_data (_T_596),	// matmul/matmul-hw.mlir:19504:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2298)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3554 (	// matmul/matmul-hw.mlir:19437:36
    .p0_rd_en   (_T_588),	// matmul/matmul-hw.mlir:19546:13
    .p1_wr_en   (_T_592),	// matmul/matmul-hw.mlir:19533:13
    .p1_wr_data (_T_591),	// matmul/matmul-hw.mlir:19534:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2297)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3555 (	// matmul/matmul-hw.mlir:19438:36
    .p0_rd_en   (_T_583),	// matmul/matmul-hw.mlir:19576:13
    .p1_wr_en   (_T_587),	// matmul/matmul-hw.mlir:19563:13
    .p1_wr_data (_T_586),	// matmul/matmul-hw.mlir:19564:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2296)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3556 (	// matmul/matmul-hw.mlir:19439:36
    .p0_rd_en   (_T_578),	// matmul/matmul-hw.mlir:19606:13
    .p1_wr_en   (_T_582),	// matmul/matmul-hw.mlir:19593:13
    .p1_wr_data (_T_581),	// matmul/matmul-hw.mlir:19594:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2295)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3557 (	// matmul/matmul-hw.mlir:19440:36
    .p0_rd_en   (_T_573),	// matmul/matmul-hw.mlir:19636:13
    .p1_wr_en   (_T_577),	// matmul/matmul-hw.mlir:19623:13
    .p1_wr_data (_T_576),	// matmul/matmul-hw.mlir:19624:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2294)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3558 (	// matmul/matmul-hw.mlir:19441:36
    .p0_rd_en   (_T_568),	// matmul/matmul-hw.mlir:19666:13
    .p1_wr_en   (_T_572),	// matmul/matmul-hw.mlir:19653:13
    .p1_wr_data (_T_571),	// matmul/matmul-hw.mlir:19654:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2293)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3559 (	// matmul/matmul-hw.mlir:19442:36
    .p0_rd_en   (_T_563),	// matmul/matmul-hw.mlir:19696:13
    .p1_wr_en   (_T_567),	// matmul/matmul-hw.mlir:19683:13
    .p1_wr_data (_T_566),	// matmul/matmul-hw.mlir:19684:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2292)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3560 (	// matmul/matmul-hw.mlir:19443:36
    .p0_rd_en   (_T_558),	// matmul/matmul-hw.mlir:19726:13
    .p1_wr_en   (_T_562),	// matmul/matmul-hw.mlir:19713:13
    .p1_wr_data (_T_561),	// matmul/matmul-hw.mlir:19714:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2291)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3561 (	// matmul/matmul-hw.mlir:19444:37
    .p0_rd_en   (_T_553),	// matmul/matmul-hw.mlir:19756:13
    .p1_wr_en   (_T_557),	// matmul/matmul-hw.mlir:19743:13
    .p1_wr_data (_T_556),	// matmul/matmul-hw.mlir:19744:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2290)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3562 (	// matmul/matmul-hw.mlir:19445:37
    .p0_rd_en   (_T_548),	// matmul/matmul-hw.mlir:19786:13
    .p1_wr_en   (_T_552),	// matmul/matmul-hw.mlir:19773:13
    .p1_wr_data (_T_551),	// matmul/matmul-hw.mlir:19774:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2289)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3563 (	// matmul/matmul-hw.mlir:19446:37
    .p0_rd_en   (_T_543),	// matmul/matmul-hw.mlir:19816:13
    .p1_wr_en   (_T_547),	// matmul/matmul-hw.mlir:19803:13
    .p1_wr_data (_T_546),	// matmul/matmul-hw.mlir:19804:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2288)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3564 (	// matmul/matmul-hw.mlir:19447:37
    .p0_rd_en   (_T_538),	// matmul/matmul-hw.mlir:19846:13
    .p1_wr_en   (_T_542),	// matmul/matmul-hw.mlir:19833:13
    .p1_wr_data (_T_541),	// matmul/matmul-hw.mlir:19834:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2287)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3565 (	// matmul/matmul-hw.mlir:19448:37
    .p0_rd_en   (_T_533),	// matmul/matmul-hw.mlir:19876:13
    .p1_wr_en   (_T_537),	// matmul/matmul-hw.mlir:19863:13
    .p1_wr_data (_T_536),	// matmul/matmul-hw.mlir:19864:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2286)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3566 (	// matmul/matmul-hw.mlir:19449:37
    .p0_rd_en   (_T_528),	// matmul/matmul-hw.mlir:19906:13
    .p1_wr_en   (_T_532),	// matmul/matmul-hw.mlir:19893:13
    .p1_wr_data (_T_531),	// matmul/matmul-hw.mlir:19894:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2285)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3567 (	// matmul/matmul-hw.mlir:19450:37
    .p0_rd_en   (_T_525),	// matmul/matmul-hw.mlir:19933:13
    .p1_wr_en   (_T_527),	// matmul/matmul-hw.mlir:19923:13
    .p1_wr_data (_T_526),	// matmul/matmul-hw.mlir:19924:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2284)
  );
  assign _T_607 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19451:13
  assign _T_606 = _T_2841 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8641:18, :19452:13
  assign _T_605 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19453:13
  assign _T_604 = _T_2830 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19454:13
  mult mult_inst144 (	// matmul/matmul-hw.mlir:19455:28
    .a      (A_reg_bank144_p0_rd_data),	// matmul/matmul-hw.mlir:12359:33
    .b      (_T_2463),
    .t      (_T_2830),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst144_result)
  );
  assign _T_603 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19456:13
  assign a_i_k_0_i_j_9 = A_reg_bank144_p0_rd_data;	// matmul/matmul-hw.mlir:12359:33, :19458:5
  //PROBE: a_i_k_0_i_j_9	// matmul/matmul-hw.mlir:19459:5
  assign b_i_k_0_i_j_9 = _T_2463;	// matmul/matmul-hw.mlir:19461:5
  //PROBE: b_i_k_0_i_j_9	// matmul/matmul-hw.mlir:19462:5
  assign c_prev_i_k_0_i_j_9 = C_reg_bank0_p0_rd_data_2300;	// matmul/matmul-hw.mlir:19434:36, :19464:5
  //PROBE: c_prev_i_k_0_i_j_9	// matmul/matmul-hw.mlir:19465:5
  assign tk_i_k_0_i_j_9 = _T_2808;	// matmul/matmul-hw.mlir:19467:5
  //PROBE: tk_i_k_0_i_j_9	// matmul/matmul-hw.mlir:19468:5
  wire [31:0] _T_3568 = mult_inst144_result + C_reg_bank0_p0_rd_data_2300;	// matmul/matmul-hw.mlir:19434:36, :19455:28, :19469:13
  assign c_i_k_0_i_j_9 = _T_3568;	// matmul/matmul-hw.mlir:19471:5
  //PROBE: c_i_k_0_i_j_9	// matmul/matmul-hw.mlir:19472:5
  assign _T_602 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19473:13
  assign _T_601 = _T_2852 ? _T_3568 : 32'bx;	// matmul/matmul-hw.mlir:8636:18, :19474:13
  localparam [3:0] _T_3570 = 4'h0;	// matmul/matmul-hw.mlir:19477:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19478:5
    if (rst)	// matmul/matmul-hw.mlir:19478:5
      i_k_next_3569 <= _T_3570;	// matmul/matmul-hw.mlir:19481:7
    else	// matmul/matmul-hw.mlir:19478:5
      i_k_next_3569 <= i_j_next_3549;	// matmul/matmul-hw.mlir:19359:13, :19479:7
  end // always @(posedge)
  assign _T_600 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19483:13
  assign _T_599 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19484:13
  mult mult_inst145 (	// matmul/matmul-hw.mlir:19485:28
    .a      (A_reg_bank145_p0_rd_data),	// matmul/matmul-hw.mlir:12360:33
    .b      (_T_2479),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst145_result)
  );
  assign _T_598 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19486:13
  assign a_i_k_1_i_j_9 = A_reg_bank145_p0_rd_data;	// matmul/matmul-hw.mlir:12360:33, :19488:5
  //PROBE: a_i_k_1_i_j_9	// matmul/matmul-hw.mlir:19489:5
  assign b_i_k_1_i_j_9 = _T_2479;	// matmul/matmul-hw.mlir:19491:5
  //PROBE: b_i_k_1_i_j_9	// matmul/matmul-hw.mlir:19492:5
  assign c_prev_i_k_1_i_j_9 = C_reg_bank1_p0_rd_data_2299;	// matmul/matmul-hw.mlir:19435:36, :19494:5
  //PROBE: c_prev_i_k_1_i_j_9	// matmul/matmul-hw.mlir:19495:5
  assign tk_i_k_1_i_j_9 = _T_2819;	// matmul/matmul-hw.mlir:19497:5
  //PROBE: tk_i_k_1_i_j_9	// matmul/matmul-hw.mlir:19498:5
  wire [31:0] _T_3571 = mult_inst145_result + C_reg_bank1_p0_rd_data_2299;	// matmul/matmul-hw.mlir:19435:36, :19485:28, :19499:13
  assign c_i_k_1_i_j_9 = _T_3571;	// matmul/matmul-hw.mlir:19501:5
  //PROBE: c_i_k_1_i_j_9	// matmul/matmul-hw.mlir:19502:5
  assign _T_597 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19503:13
  assign _T_596 = _T_2863 ? _T_3571 : 32'bx;	// matmul/matmul-hw.mlir:8631:18, :19504:13
  localparam [3:0] _T_3573 = 4'h0;	// matmul/matmul-hw.mlir:19507:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19508:5
    if (rst)	// matmul/matmul-hw.mlir:19508:5
      i_k_next_3572 <= _T_3573;	// matmul/matmul-hw.mlir:19511:7
    else	// matmul/matmul-hw.mlir:19508:5
      i_k_next_3572 <= i_k_next_3569;	// matmul/matmul-hw.mlir:19476:13, :19509:7
  end // always @(posedge)
  assign _T_595 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19513:13
  assign _T_594 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19514:13
  mult mult_inst146 (	// matmul/matmul-hw.mlir:19515:28
    .a      (A_reg_bank146_p0_rd_data),	// matmul/matmul-hw.mlir:12361:33
    .b      (_T_2495),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst146_result)
  );
  assign _T_593 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19516:13
  assign a_i_k_2_i_j_9 = A_reg_bank146_p0_rd_data;	// matmul/matmul-hw.mlir:12361:33, :19518:5
  //PROBE: a_i_k_2_i_j_9	// matmul/matmul-hw.mlir:19519:5
  assign b_i_k_2_i_j_9 = _T_2495;	// matmul/matmul-hw.mlir:19521:5
  //PROBE: b_i_k_2_i_j_9	// matmul/matmul-hw.mlir:19522:5
  assign c_prev_i_k_2_i_j_9 = C_reg_bank2_p0_rd_data_2298;	// matmul/matmul-hw.mlir:19436:36, :19524:5
  //PROBE: c_prev_i_k_2_i_j_9	// matmul/matmul-hw.mlir:19525:5
  assign tk_i_k_2_i_j_9 = _T_2830;	// matmul/matmul-hw.mlir:19527:5
  //PROBE: tk_i_k_2_i_j_9	// matmul/matmul-hw.mlir:19528:5
  wire [31:0] _T_3574 = mult_inst146_result + C_reg_bank2_p0_rd_data_2298;	// matmul/matmul-hw.mlir:19436:36, :19515:28, :19529:13
  assign c_i_k_2_i_j_9 = _T_3574;	// matmul/matmul-hw.mlir:19531:5
  //PROBE: c_i_k_2_i_j_9	// matmul/matmul-hw.mlir:19532:5
  assign _T_592 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19533:13
  assign _T_591 = _T_2874 ? _T_3574 : 32'bx;	// matmul/matmul-hw.mlir:8626:18, :19534:13
  localparam [3:0] _T_3576 = 4'h0;	// matmul/matmul-hw.mlir:19537:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19538:5
    if (rst)	// matmul/matmul-hw.mlir:19538:5
      i_k_next_3575 <= _T_3576;	// matmul/matmul-hw.mlir:19541:7
    else	// matmul/matmul-hw.mlir:19538:5
      i_k_next_3575 <= i_k_next_3572;	// matmul/matmul-hw.mlir:19506:13, :19539:7
  end // always @(posedge)
  assign _T_590 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19543:13
  assign _T_589 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19544:13
  mult mult_inst147 (	// matmul/matmul-hw.mlir:19545:28
    .a      (A_reg_bank147_p0_rd_data),	// matmul/matmul-hw.mlir:12362:33
    .b      (_T_2511),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst147_result)
  );
  assign _T_588 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19546:13
  assign a_i_k_3_i_j_9 = A_reg_bank147_p0_rd_data;	// matmul/matmul-hw.mlir:12362:33, :19548:5
  //PROBE: a_i_k_3_i_j_9	// matmul/matmul-hw.mlir:19549:5
  assign b_i_k_3_i_j_9 = _T_2511;	// matmul/matmul-hw.mlir:19551:5
  //PROBE: b_i_k_3_i_j_9	// matmul/matmul-hw.mlir:19552:5
  assign c_prev_i_k_3_i_j_9 = C_reg_bank3_p0_rd_data_2297;	// matmul/matmul-hw.mlir:19437:36, :19554:5
  //PROBE: c_prev_i_k_3_i_j_9	// matmul/matmul-hw.mlir:19555:5
  assign tk_i_k_3_i_j_9 = _T_2841;	// matmul/matmul-hw.mlir:19557:5
  //PROBE: tk_i_k_3_i_j_9	// matmul/matmul-hw.mlir:19558:5
  wire [31:0] _T_3577 = mult_inst147_result + C_reg_bank3_p0_rd_data_2297;	// matmul/matmul-hw.mlir:19437:36, :19545:28, :19559:13
  assign c_i_k_3_i_j_9 = _T_3577;	// matmul/matmul-hw.mlir:19561:5
  //PROBE: c_i_k_3_i_j_9	// matmul/matmul-hw.mlir:19562:5
  assign _T_587 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19563:13
  assign _T_586 = _T_2885 ? _T_3577 : 32'bx;	// matmul/matmul-hw.mlir:8621:18, :19564:13
  localparam [3:0] _T_3579 = 4'h0;	// matmul/matmul-hw.mlir:19567:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19568:5
    if (rst)	// matmul/matmul-hw.mlir:19568:5
      i_k_next_3578 <= _T_3579;	// matmul/matmul-hw.mlir:19571:7
    else	// matmul/matmul-hw.mlir:19568:5
      i_k_next_3578 <= i_k_next_3575;	// matmul/matmul-hw.mlir:19536:13, :19569:7
  end // always @(posedge)
  assign _T_585 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19573:13
  assign _T_584 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19574:13
  mult mult_inst148 (	// matmul/matmul-hw.mlir:19575:28
    .a      (A_reg_bank148_p0_rd_data),	// matmul/matmul-hw.mlir:12363:33
    .b      (_T_2527),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst148_result)
  );
  assign _T_583 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19576:13
  assign a_i_k_4_i_j_9 = A_reg_bank148_p0_rd_data;	// matmul/matmul-hw.mlir:12363:33, :19578:5
  //PROBE: a_i_k_4_i_j_9	// matmul/matmul-hw.mlir:19579:5
  assign b_i_k_4_i_j_9 = _T_2527;	// matmul/matmul-hw.mlir:19581:5
  //PROBE: b_i_k_4_i_j_9	// matmul/matmul-hw.mlir:19582:5
  assign c_prev_i_k_4_i_j_9 = C_reg_bank4_p0_rd_data_2296;	// matmul/matmul-hw.mlir:19438:36, :19584:5
  //PROBE: c_prev_i_k_4_i_j_9	// matmul/matmul-hw.mlir:19585:5
  assign tk_i_k_4_i_j_9 = _T_2852;	// matmul/matmul-hw.mlir:19587:5
  //PROBE: tk_i_k_4_i_j_9	// matmul/matmul-hw.mlir:19588:5
  wire [31:0] _T_3580 = mult_inst148_result + C_reg_bank4_p0_rd_data_2296;	// matmul/matmul-hw.mlir:19438:36, :19575:28, :19589:13
  assign c_i_k_4_i_j_9 = _T_3580;	// matmul/matmul-hw.mlir:19591:5
  //PROBE: c_i_k_4_i_j_9	// matmul/matmul-hw.mlir:19592:5
  assign _T_582 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19593:13
  assign _T_581 = _T_2892 ? _T_3580 : 32'bx;	// matmul/matmul-hw.mlir:8616:18, :19594:13
  localparam [3:0] _T_3582 = 4'h0;	// matmul/matmul-hw.mlir:19597:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19598:5
    if (rst)	// matmul/matmul-hw.mlir:19598:5
      i_k_next_3581 <= _T_3582;	// matmul/matmul-hw.mlir:19601:7
    else	// matmul/matmul-hw.mlir:19598:5
      i_k_next_3581 <= i_k_next_3578;	// matmul/matmul-hw.mlir:19566:13, :19599:7
  end // always @(posedge)
  assign _T_580 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19603:13
  assign _T_579 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19604:13
  mult mult_inst149 (	// matmul/matmul-hw.mlir:19605:28
    .a      (A_reg_bank149_p0_rd_data),	// matmul/matmul-hw.mlir:12364:33
    .b      (_T_2543),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst149_result)
  );
  assign _T_578 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19606:13
  assign a_i_k_5_i_j_9 = A_reg_bank149_p0_rd_data;	// matmul/matmul-hw.mlir:12364:33, :19608:5
  //PROBE: a_i_k_5_i_j_9	// matmul/matmul-hw.mlir:19609:5
  assign b_i_k_5_i_j_9 = _T_2543;	// matmul/matmul-hw.mlir:19611:5
  //PROBE: b_i_k_5_i_j_9	// matmul/matmul-hw.mlir:19612:5
  assign c_prev_i_k_5_i_j_9 = C_reg_bank5_p0_rd_data_2295;	// matmul/matmul-hw.mlir:19439:36, :19614:5
  //PROBE: c_prev_i_k_5_i_j_9	// matmul/matmul-hw.mlir:19615:5
  assign tk_i_k_5_i_j_9 = _T_2863;	// matmul/matmul-hw.mlir:19617:5
  //PROBE: tk_i_k_5_i_j_9	// matmul/matmul-hw.mlir:19618:5
  wire [31:0] _T_3583 = mult_inst149_result + C_reg_bank5_p0_rd_data_2295;	// matmul/matmul-hw.mlir:19439:36, :19605:28, :19619:13
  assign c_i_k_5_i_j_9 = _T_3583;	// matmul/matmul-hw.mlir:19621:5
  //PROBE: c_i_k_5_i_j_9	// matmul/matmul-hw.mlir:19622:5
  assign _T_577 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19623:13
  assign _T_576 = _T_2897 ? _T_3583 : 32'bx;	// matmul/matmul-hw.mlir:8611:18, :19624:13
  localparam [3:0] _T_3585 = 4'h0;	// matmul/matmul-hw.mlir:19627:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19628:5
    if (rst)	// matmul/matmul-hw.mlir:19628:5
      i_k_next_3584 <= _T_3585;	// matmul/matmul-hw.mlir:19631:7
    else	// matmul/matmul-hw.mlir:19628:5
      i_k_next_3584 <= i_k_next_3581;	// matmul/matmul-hw.mlir:19596:13, :19629:7
  end // always @(posedge)
  assign _T_575 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19633:13
  assign _T_574 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19634:13
  mult mult_inst150 (	// matmul/matmul-hw.mlir:19635:28
    .a      (A_reg_bank150_p0_rd_data),	// matmul/matmul-hw.mlir:12365:33
    .b      (_T_2559),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst150_result)
  );
  assign _T_573 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19636:13
  assign a_i_k_6_i_j_9 = A_reg_bank150_p0_rd_data;	// matmul/matmul-hw.mlir:12365:33, :19638:5
  //PROBE: a_i_k_6_i_j_9	// matmul/matmul-hw.mlir:19639:5
  assign b_i_k_6_i_j_9 = _T_2559;	// matmul/matmul-hw.mlir:19641:5
  //PROBE: b_i_k_6_i_j_9	// matmul/matmul-hw.mlir:19642:5
  assign c_prev_i_k_6_i_j_9 = C_reg_bank6_p0_rd_data_2294;	// matmul/matmul-hw.mlir:19440:36, :19644:5
  //PROBE: c_prev_i_k_6_i_j_9	// matmul/matmul-hw.mlir:19645:5
  assign tk_i_k_6_i_j_9 = _T_2874;	// matmul/matmul-hw.mlir:19647:5
  //PROBE: tk_i_k_6_i_j_9	// matmul/matmul-hw.mlir:19648:5
  wire [31:0] _T_3586 = mult_inst150_result + C_reg_bank6_p0_rd_data_2294;	// matmul/matmul-hw.mlir:19440:36, :19635:28, :19649:13
  assign c_i_k_6_i_j_9 = _T_3586;	// matmul/matmul-hw.mlir:19651:5
  //PROBE: c_i_k_6_i_j_9	// matmul/matmul-hw.mlir:19652:5
  assign _T_572 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19653:13
  assign _T_571 = _T_2902 ? _T_3586 : 32'bx;	// matmul/matmul-hw.mlir:8606:18, :19654:13
  localparam [3:0] _T_3588 = 4'h0;	// matmul/matmul-hw.mlir:19657:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19658:5
    if (rst)	// matmul/matmul-hw.mlir:19658:5
      i_k_next_3587 <= _T_3588;	// matmul/matmul-hw.mlir:19661:7
    else	// matmul/matmul-hw.mlir:19658:5
      i_k_next_3587 <= i_k_next_3584;	// matmul/matmul-hw.mlir:19626:13, :19659:7
  end // always @(posedge)
  assign _T_570 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19663:13
  assign _T_569 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19664:13
  mult mult_inst151 (	// matmul/matmul-hw.mlir:19665:28
    .a      (A_reg_bank151_p0_rd_data),	// matmul/matmul-hw.mlir:12366:33
    .b      (_T_2575),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst151_result)
  );
  assign _T_568 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19666:13
  assign a_i_k_7_i_j_9 = A_reg_bank151_p0_rd_data;	// matmul/matmul-hw.mlir:12366:33, :19668:5
  //PROBE: a_i_k_7_i_j_9	// matmul/matmul-hw.mlir:19669:5
  assign b_i_k_7_i_j_9 = _T_2575;	// matmul/matmul-hw.mlir:19671:5
  //PROBE: b_i_k_7_i_j_9	// matmul/matmul-hw.mlir:19672:5
  assign c_prev_i_k_7_i_j_9 = C_reg_bank7_p0_rd_data_2293;	// matmul/matmul-hw.mlir:19441:36, :19674:5
  //PROBE: c_prev_i_k_7_i_j_9	// matmul/matmul-hw.mlir:19675:5
  assign tk_i_k_7_i_j_9 = _T_2885;	// matmul/matmul-hw.mlir:19677:5
  //PROBE: tk_i_k_7_i_j_9	// matmul/matmul-hw.mlir:19678:5
  wire [31:0] _T_3589 = mult_inst151_result + C_reg_bank7_p0_rd_data_2293;	// matmul/matmul-hw.mlir:19441:36, :19665:28, :19679:13
  assign c_i_k_7_i_j_9 = _T_3589;	// matmul/matmul-hw.mlir:19681:5
  //PROBE: c_i_k_7_i_j_9	// matmul/matmul-hw.mlir:19682:5
  assign _T_567 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19683:13
  assign _T_566 = _T_2907 ? _T_3589 : 32'bx;	// matmul/matmul-hw.mlir:8601:18, :19684:13
  localparam [3:0] _T_3591 = 4'h0;	// matmul/matmul-hw.mlir:19687:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19688:5
    if (rst)	// matmul/matmul-hw.mlir:19688:5
      i_k_next_3590 <= _T_3591;	// matmul/matmul-hw.mlir:19691:7
    else	// matmul/matmul-hw.mlir:19688:5
      i_k_next_3590 <= i_k_next_3587;	// matmul/matmul-hw.mlir:19656:13, :19689:7
  end // always @(posedge)
  assign _T_565 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19693:13
  assign _T_564 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19694:13
  mult mult_inst152 (	// matmul/matmul-hw.mlir:19695:28
    .a      (A_reg_bank152_p0_rd_data),	// matmul/matmul-hw.mlir:12367:33
    .b      (_T_2591),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst152_result)
  );
  assign _T_563 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19696:13
  assign a_i_k_8_i_j_9 = A_reg_bank152_p0_rd_data;	// matmul/matmul-hw.mlir:12367:33, :19698:5
  //PROBE: a_i_k_8_i_j_9	// matmul/matmul-hw.mlir:19699:5
  assign b_i_k_8_i_j_9 = _T_2591;	// matmul/matmul-hw.mlir:19701:5
  //PROBE: b_i_k_8_i_j_9	// matmul/matmul-hw.mlir:19702:5
  assign c_prev_i_k_8_i_j_9 = C_reg_bank8_p0_rd_data_2292;	// matmul/matmul-hw.mlir:19442:36, :19704:5
  //PROBE: c_prev_i_k_8_i_j_9	// matmul/matmul-hw.mlir:19705:5
  assign tk_i_k_8_i_j_9 = _T_2892;	// matmul/matmul-hw.mlir:19707:5
  //PROBE: tk_i_k_8_i_j_9	// matmul/matmul-hw.mlir:19708:5
  wire [31:0] _T_3592 = mult_inst152_result + C_reg_bank8_p0_rd_data_2292;	// matmul/matmul-hw.mlir:19442:36, :19695:28, :19709:13
  assign c_i_k_8_i_j_9 = _T_3592;	// matmul/matmul-hw.mlir:19711:5
  //PROBE: c_i_k_8_i_j_9	// matmul/matmul-hw.mlir:19712:5
  assign _T_562 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19713:13
  assign _T_561 = _T_2912 ? _T_3592 : 32'bx;	// matmul/matmul-hw.mlir:8596:18, :19714:13
  localparam [3:0] _T_3594 = 4'h0;	// matmul/matmul-hw.mlir:19717:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19718:5
    if (rst)	// matmul/matmul-hw.mlir:19718:5
      i_k_next_3593 <= _T_3594;	// matmul/matmul-hw.mlir:19721:7
    else	// matmul/matmul-hw.mlir:19718:5
      i_k_next_3593 <= i_k_next_3590;	// matmul/matmul-hw.mlir:19686:13, :19719:7
  end // always @(posedge)
  assign _T_560 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19723:13
  assign _T_559 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19724:13
  mult mult_inst153 (	// matmul/matmul-hw.mlir:19725:28
    .a      (A_reg_bank153_p0_rd_data),	// matmul/matmul-hw.mlir:12368:33
    .b      (_T_2607),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst153_result)
  );
  assign _T_558 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19726:13
  assign a_i_k_9_i_j_9 = A_reg_bank153_p0_rd_data;	// matmul/matmul-hw.mlir:12368:33, :19728:5
  //PROBE: a_i_k_9_i_j_9	// matmul/matmul-hw.mlir:19729:5
  assign b_i_k_9_i_j_9 = _T_2607;	// matmul/matmul-hw.mlir:19731:5
  //PROBE: b_i_k_9_i_j_9	// matmul/matmul-hw.mlir:19732:5
  assign c_prev_i_k_9_i_j_9 = C_reg_bank9_p0_rd_data_2291;	// matmul/matmul-hw.mlir:19443:36, :19734:5
  //PROBE: c_prev_i_k_9_i_j_9	// matmul/matmul-hw.mlir:19735:5
  assign tk_i_k_9_i_j_9 = _T_2897;	// matmul/matmul-hw.mlir:19737:5
  //PROBE: tk_i_k_9_i_j_9	// matmul/matmul-hw.mlir:19738:5
  wire [31:0] _T_3595 = mult_inst153_result + C_reg_bank9_p0_rd_data_2291;	// matmul/matmul-hw.mlir:19443:36, :19725:28, :19739:13
  assign c_i_k_9_i_j_9 = _T_3595;	// matmul/matmul-hw.mlir:19741:5
  //PROBE: c_i_k_9_i_j_9	// matmul/matmul-hw.mlir:19742:5
  assign _T_557 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19743:13
  assign _T_556 = _T_2917 ? _T_3595 : 32'bx;	// matmul/matmul-hw.mlir:8591:18, :19744:13
  localparam [3:0] _T_3597 = 4'h0;	// matmul/matmul-hw.mlir:19747:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19748:5
    if (rst)	// matmul/matmul-hw.mlir:19748:5
      i_k_next_3596 <= _T_3597;	// matmul/matmul-hw.mlir:19751:7
    else	// matmul/matmul-hw.mlir:19748:5
      i_k_next_3596 <= i_k_next_3593;	// matmul/matmul-hw.mlir:19716:13, :19749:7
  end // always @(posedge)
  assign _T_555 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19753:13
  assign _T_554 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19754:13
  mult mult_inst154 (	// matmul/matmul-hw.mlir:19755:28
    .a      (A_reg_bank154_p0_rd_data),	// matmul/matmul-hw.mlir:12369:33
    .b      (_T_2623),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst154_result)
  );
  assign _T_553 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19756:13
  assign a_i_k_10_i_j_9 = A_reg_bank154_p0_rd_data;	// matmul/matmul-hw.mlir:12369:33, :19758:5
  //PROBE: a_i_k_10_i_j_9	// matmul/matmul-hw.mlir:19759:5
  assign b_i_k_10_i_j_9 = _T_2623;	// matmul/matmul-hw.mlir:19761:5
  //PROBE: b_i_k_10_i_j_9	// matmul/matmul-hw.mlir:19762:5
  assign c_prev_i_k_10_i_j_9 = C_reg_bank10_p0_rd_data_2290;	// matmul/matmul-hw.mlir:19444:37, :19764:5
  //PROBE: c_prev_i_k_10_i_j_9	// matmul/matmul-hw.mlir:19765:5
  assign tk_i_k_10_i_j_9 = _T_2902;	// matmul/matmul-hw.mlir:19767:5
  //PROBE: tk_i_k_10_i_j_9	// matmul/matmul-hw.mlir:19768:5
  wire [31:0] _T_3598 = mult_inst154_result + C_reg_bank10_p0_rd_data_2290;	// matmul/matmul-hw.mlir:19444:37, :19755:28, :19769:13
  assign c_i_k_10_i_j_9 = _T_3598;	// matmul/matmul-hw.mlir:19771:5
  //PROBE: c_i_k_10_i_j_9	// matmul/matmul-hw.mlir:19772:5
  assign _T_552 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19773:13
  assign _T_551 = _T_2922 ? _T_3598 : 32'bx;	// matmul/matmul-hw.mlir:8586:18, :19774:13
  localparam [3:0] _T_3600 = 4'h0;	// matmul/matmul-hw.mlir:19777:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19778:5
    if (rst)	// matmul/matmul-hw.mlir:19778:5
      i_k_next_3599 <= _T_3600;	// matmul/matmul-hw.mlir:19781:7
    else	// matmul/matmul-hw.mlir:19778:5
      i_k_next_3599 <= i_k_next_3596;	// matmul/matmul-hw.mlir:19746:13, :19779:7
  end // always @(posedge)
  assign _T_550 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19783:13
  assign _T_549 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19784:13
  mult mult_inst155 (	// matmul/matmul-hw.mlir:19785:28
    .a      (A_reg_bank155_p0_rd_data),	// matmul/matmul-hw.mlir:12370:33
    .b      (_T_2639),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst155_result)
  );
  assign _T_548 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19786:13
  assign a_i_k_11_i_j_9 = A_reg_bank155_p0_rd_data;	// matmul/matmul-hw.mlir:12370:33, :19788:5
  //PROBE: a_i_k_11_i_j_9	// matmul/matmul-hw.mlir:19789:5
  assign b_i_k_11_i_j_9 = _T_2639;	// matmul/matmul-hw.mlir:19791:5
  //PROBE: b_i_k_11_i_j_9	// matmul/matmul-hw.mlir:19792:5
  assign c_prev_i_k_11_i_j_9 = C_reg_bank11_p0_rd_data_2289;	// matmul/matmul-hw.mlir:19445:37, :19794:5
  //PROBE: c_prev_i_k_11_i_j_9	// matmul/matmul-hw.mlir:19795:5
  assign tk_i_k_11_i_j_9 = _T_2907;	// matmul/matmul-hw.mlir:19797:5
  //PROBE: tk_i_k_11_i_j_9	// matmul/matmul-hw.mlir:19798:5
  wire [31:0] _T_3601 = mult_inst155_result + C_reg_bank11_p0_rd_data_2289;	// matmul/matmul-hw.mlir:19445:37, :19785:28, :19799:13
  assign c_i_k_11_i_j_9 = _T_3601;	// matmul/matmul-hw.mlir:19801:5
  //PROBE: c_i_k_11_i_j_9	// matmul/matmul-hw.mlir:19802:5
  assign _T_547 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19803:13
  assign _T_546 = _T_2927 ? _T_3601 : 32'bx;	// matmul/matmul-hw.mlir:8581:18, :19804:13
  localparam [3:0] _T_3603 = 4'h0;	// matmul/matmul-hw.mlir:19807:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19808:5
    if (rst)	// matmul/matmul-hw.mlir:19808:5
      i_k_next_3602 <= _T_3603;	// matmul/matmul-hw.mlir:19811:7
    else	// matmul/matmul-hw.mlir:19808:5
      i_k_next_3602 <= i_k_next_3599;	// matmul/matmul-hw.mlir:19776:13, :19809:7
  end // always @(posedge)
  assign _T_545 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19813:13
  assign _T_544 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19814:13
  mult mult_inst156 (	// matmul/matmul-hw.mlir:19815:28
    .a      (A_reg_bank156_p0_rd_data),	// matmul/matmul-hw.mlir:12371:33
    .b      (_T_2655),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst156_result)
  );
  assign _T_543 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19816:13
  assign a_i_k_12_i_j_9 = A_reg_bank156_p0_rd_data;	// matmul/matmul-hw.mlir:12371:33, :19818:5
  //PROBE: a_i_k_12_i_j_9	// matmul/matmul-hw.mlir:19819:5
  assign b_i_k_12_i_j_9 = _T_2655;	// matmul/matmul-hw.mlir:19821:5
  //PROBE: b_i_k_12_i_j_9	// matmul/matmul-hw.mlir:19822:5
  assign c_prev_i_k_12_i_j_9 = C_reg_bank12_p0_rd_data_2288;	// matmul/matmul-hw.mlir:19446:37, :19824:5
  //PROBE: c_prev_i_k_12_i_j_9	// matmul/matmul-hw.mlir:19825:5
  assign tk_i_k_12_i_j_9 = _T_2912;	// matmul/matmul-hw.mlir:19827:5
  //PROBE: tk_i_k_12_i_j_9	// matmul/matmul-hw.mlir:19828:5
  wire [31:0] _T_3604 = mult_inst156_result + C_reg_bank12_p0_rd_data_2288;	// matmul/matmul-hw.mlir:19446:37, :19815:28, :19829:13
  assign c_i_k_12_i_j_9 = _T_3604;	// matmul/matmul-hw.mlir:19831:5
  //PROBE: c_i_k_12_i_j_9	// matmul/matmul-hw.mlir:19832:5
  assign _T_542 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19833:13
  assign _T_541 = _T_2932 ? _T_3604 : 32'bx;	// matmul/matmul-hw.mlir:8576:18, :19834:13
  localparam [3:0] _T_3606 = 4'h0;	// matmul/matmul-hw.mlir:19837:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19838:5
    if (rst)	// matmul/matmul-hw.mlir:19838:5
      i_k_next_3605 <= _T_3606;	// matmul/matmul-hw.mlir:19841:7
    else	// matmul/matmul-hw.mlir:19838:5
      i_k_next_3605 <= i_k_next_3602;	// matmul/matmul-hw.mlir:19806:13, :19839:7
  end // always @(posedge)
  assign _T_540 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19843:13
  assign _T_539 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19844:13
  mult mult_inst157 (	// matmul/matmul-hw.mlir:19845:28
    .a      (A_reg_bank157_p0_rd_data),	// matmul/matmul-hw.mlir:12372:33
    .b      (_T_2671),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst157_result)
  );
  assign _T_538 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19846:13
  assign a_i_k_13_i_j_9 = A_reg_bank157_p0_rd_data;	// matmul/matmul-hw.mlir:12372:33, :19848:5
  //PROBE: a_i_k_13_i_j_9	// matmul/matmul-hw.mlir:19849:5
  assign b_i_k_13_i_j_9 = _T_2671;	// matmul/matmul-hw.mlir:19851:5
  //PROBE: b_i_k_13_i_j_9	// matmul/matmul-hw.mlir:19852:5
  assign c_prev_i_k_13_i_j_9 = C_reg_bank13_p0_rd_data_2287;	// matmul/matmul-hw.mlir:19447:37, :19854:5
  //PROBE: c_prev_i_k_13_i_j_9	// matmul/matmul-hw.mlir:19855:5
  assign tk_i_k_13_i_j_9 = _T_2917;	// matmul/matmul-hw.mlir:19857:5
  //PROBE: tk_i_k_13_i_j_9	// matmul/matmul-hw.mlir:19858:5
  wire [31:0] _T_3607 = mult_inst157_result + C_reg_bank13_p0_rd_data_2287;	// matmul/matmul-hw.mlir:19447:37, :19845:28, :19859:13
  assign c_i_k_13_i_j_9 = _T_3607;	// matmul/matmul-hw.mlir:19861:5
  //PROBE: c_i_k_13_i_j_9	// matmul/matmul-hw.mlir:19862:5
  assign _T_537 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19863:13
  assign _T_536 = _T_2937 ? _T_3607 : 32'bx;	// matmul/matmul-hw.mlir:8571:18, :19864:13
  localparam [3:0] _T_3609 = 4'h0;	// matmul/matmul-hw.mlir:19867:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19868:5
    if (rst)	// matmul/matmul-hw.mlir:19868:5
      i_k_next_3608 <= _T_3609;	// matmul/matmul-hw.mlir:19871:7
    else	// matmul/matmul-hw.mlir:19868:5
      i_k_next_3608 <= i_k_next_3605;	// matmul/matmul-hw.mlir:19836:13, :19869:7
  end // always @(posedge)
  assign _T_535 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19873:13
  assign _T_534 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19874:13
  mult mult_inst158 (	// matmul/matmul-hw.mlir:19875:28
    .a      (A_reg_bank158_p0_rd_data),	// matmul/matmul-hw.mlir:12373:33
    .b      (_T_2687),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst158_result)
  );
  assign _T_533 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19876:13
  assign a_i_k_14_i_j_9 = A_reg_bank158_p0_rd_data;	// matmul/matmul-hw.mlir:12373:33, :19878:5
  //PROBE: a_i_k_14_i_j_9	// matmul/matmul-hw.mlir:19879:5
  assign b_i_k_14_i_j_9 = _T_2687;	// matmul/matmul-hw.mlir:19881:5
  //PROBE: b_i_k_14_i_j_9	// matmul/matmul-hw.mlir:19882:5
  assign c_prev_i_k_14_i_j_9 = C_reg_bank14_p0_rd_data_2286;	// matmul/matmul-hw.mlir:19448:37, :19884:5
  //PROBE: c_prev_i_k_14_i_j_9	// matmul/matmul-hw.mlir:19885:5
  assign tk_i_k_14_i_j_9 = _T_2922;	// matmul/matmul-hw.mlir:19887:5
  //PROBE: tk_i_k_14_i_j_9	// matmul/matmul-hw.mlir:19888:5
  wire [31:0] _T_3610 = mult_inst158_result + C_reg_bank14_p0_rd_data_2286;	// matmul/matmul-hw.mlir:19448:37, :19875:28, :19889:13
  assign c_i_k_14_i_j_9 = _T_3610;	// matmul/matmul-hw.mlir:19891:5
  //PROBE: c_i_k_14_i_j_9	// matmul/matmul-hw.mlir:19892:5
  assign _T_532 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19893:13
  assign _T_531 = _T_2942 ? _T_3610 : 32'bx;	// matmul/matmul-hw.mlir:8566:18, :19894:13
  localparam [3:0] _T_3612 = 4'h0;	// matmul/matmul-hw.mlir:19897:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19898:5
    if (rst)	// matmul/matmul-hw.mlir:19898:5
      i_k_next_3611 <= _T_3612;	// matmul/matmul-hw.mlir:19901:7
    else	// matmul/matmul-hw.mlir:19898:5
      i_k_next_3611 <= i_k_next_3608;	// matmul/matmul-hw.mlir:19866:13, :19899:7
  end // always @(posedge)
  assign _T_530 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19903:13
  assign _T_529 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19904:13
  mult mult_inst159 (	// matmul/matmul-hw.mlir:19905:28
    .a      (A_reg_bank159_p0_rd_data),	// matmul/matmul-hw.mlir:12374:33
    .b      (_T_2703),
    .t      (_T_2937),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst159_result)
  );
  assign _T_528 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19906:13
  assign a_i_k_15_i_j_9 = A_reg_bank159_p0_rd_data;	// matmul/matmul-hw.mlir:12374:33, :19908:5
  //PROBE: a_i_k_15_i_j_9	// matmul/matmul-hw.mlir:19909:5
  assign b_i_k_15_i_j_9 = _T_2703;	// matmul/matmul-hw.mlir:19911:5
  //PROBE: b_i_k_15_i_j_9	// matmul/matmul-hw.mlir:19912:5
  assign c_prev_i_k_15_i_j_9 = C_reg_bank15_p0_rd_data_2285;	// matmul/matmul-hw.mlir:19449:37, :19914:5
  //PROBE: c_prev_i_k_15_i_j_9	// matmul/matmul-hw.mlir:19915:5
  assign tk_i_k_15_i_j_9 = _T_2927;	// matmul/matmul-hw.mlir:19917:5
  //PROBE: tk_i_k_15_i_j_9	// matmul/matmul-hw.mlir:19918:5
  wire [31:0] _T_3613 = mult_inst159_result + C_reg_bank15_p0_rd_data_2285;	// matmul/matmul-hw.mlir:19449:37, :19905:28, :19919:13
  assign c_i_k_15_i_j_9 = _T_3613;	// matmul/matmul-hw.mlir:19921:5
  //PROBE: c_i_k_15_i_j_9	// matmul/matmul-hw.mlir:19922:5
  assign _T_527 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19923:13
  assign _T_526 = _T_2947 ? _T_3613 : 32'bx;	// matmul/matmul-hw.mlir:8561:18, :19924:13
  localparam [3:0] _T_3615 = 4'h0;	// matmul/matmul-hw.mlir:19927:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19928:5
    if (rst)	// matmul/matmul-hw.mlir:19928:5
      i_k_next_3614 <= _T_3615;	// matmul/matmul-hw.mlir:19931:7
    else	// matmul/matmul-hw.mlir:19928:5
      i_k_next_3614 <= i_k_next_3611;	// matmul/matmul-hw.mlir:19896:13, :19929:7
  end // always @(posedge)
  assign _T_525 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19933:13
  wire [3:0][3:0] _T_3617 = i_delayed_3616;	// matmul/matmul-hw.mlir:19935:13
  wire [3:0][3:0] _T_3618 = {_T_3617[2'h0+:3], {{i_k_next_3614}}};	// matmul/matmul-hw.mlir:19926:13, :19936:19, :19937:13, :19938:13, :19939:13
  wire [3:0][3:0] _T_3619 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:19940:19, :19941:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19942:5
    if (rst)	// matmul/matmul-hw.mlir:19942:5
      i_delayed_3616 <= _T_3619;	// matmul/matmul-hw.mlir:19945:7
    else	// matmul/matmul-hw.mlir:19942:5
      i_delayed_3616 <= _T_3618;	// matmul/matmul-hw.mlir:19943:7
  end // always @(posedge)
  assign _T_524 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19949:13
  assign _T_523 = _T_2952 ? i_delayed_3616[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8558:17, :19935:13, :19947:20, :19948:13, :19950:13
  assign _T_522 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :19951:13
  assign _T_521 = _T_2952 ? C_reg_bank16_p0_rd_data_2284 : 32'bx;	// matmul/matmul-hw.mlir:8556:18, :19450:37, :19952:13
  localparam [3:0] _T_3621 = 4'h0;	// matmul/matmul-hw.mlir:19955:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:19956:5
    if (rst)	// matmul/matmul-hw.mlir:19956:5
      i_j_next_3620 <= _T_3621;	// matmul/matmul-hw.mlir:19959:7
    else	// matmul/matmul-hw.mlir:19956:5
      i_j_next_3620 <= i_j_next_3549;	// matmul/matmul-hw.mlir:19359:13, :19957:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3622 (	// matmul/matmul-hw.mlir:20029:36
    .p0_rd_en   (_T_516),	// matmul/matmul-hw.mlir:20051:13
    .p1_wr_en   (_T_520),	// matmul/matmul-hw.mlir:20046:13
    .p1_wr_data (_T_519),	// matmul/matmul-hw.mlir:20047:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2283)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3623 (	// matmul/matmul-hw.mlir:20030:36
    .p0_rd_en   (_T_511),	// matmul/matmul-hw.mlir:20081:13
    .p1_wr_en   (_T_515),	// matmul/matmul-hw.mlir:20068:13
    .p1_wr_data (_T_514),	// matmul/matmul-hw.mlir:20069:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2282)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3624 (	// matmul/matmul-hw.mlir:20031:36
    .p0_rd_en   (_T_506),	// matmul/matmul-hw.mlir:20111:13
    .p1_wr_en   (_T_510),	// matmul/matmul-hw.mlir:20098:13
    .p1_wr_data (_T_509),	// matmul/matmul-hw.mlir:20099:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2281)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3625 (	// matmul/matmul-hw.mlir:20032:36
    .p0_rd_en   (_T_501),	// matmul/matmul-hw.mlir:20141:13
    .p1_wr_en   (_T_505),	// matmul/matmul-hw.mlir:20128:13
    .p1_wr_data (_T_504),	// matmul/matmul-hw.mlir:20129:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2280)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3626 (	// matmul/matmul-hw.mlir:20033:36
    .p0_rd_en   (_T_496),	// matmul/matmul-hw.mlir:20171:13
    .p1_wr_en   (_T_500),	// matmul/matmul-hw.mlir:20158:13
    .p1_wr_data (_T_499),	// matmul/matmul-hw.mlir:20159:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2279)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3627 (	// matmul/matmul-hw.mlir:20034:36
    .p0_rd_en   (_T_491),	// matmul/matmul-hw.mlir:20201:13
    .p1_wr_en   (_T_495),	// matmul/matmul-hw.mlir:20188:13
    .p1_wr_data (_T_494),	// matmul/matmul-hw.mlir:20189:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2278)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3628 (	// matmul/matmul-hw.mlir:20035:36
    .p0_rd_en   (_T_486),	// matmul/matmul-hw.mlir:20231:13
    .p1_wr_en   (_T_490),	// matmul/matmul-hw.mlir:20218:13
    .p1_wr_data (_T_489),	// matmul/matmul-hw.mlir:20219:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2277)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3629 (	// matmul/matmul-hw.mlir:20036:36
    .p0_rd_en   (_T_481),	// matmul/matmul-hw.mlir:20261:13
    .p1_wr_en   (_T_485),	// matmul/matmul-hw.mlir:20248:13
    .p1_wr_data (_T_484),	// matmul/matmul-hw.mlir:20249:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2276)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3630 (	// matmul/matmul-hw.mlir:20037:36
    .p0_rd_en   (_T_476),	// matmul/matmul-hw.mlir:20291:13
    .p1_wr_en   (_T_480),	// matmul/matmul-hw.mlir:20278:13
    .p1_wr_data (_T_479),	// matmul/matmul-hw.mlir:20279:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2275)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3631 (	// matmul/matmul-hw.mlir:20038:36
    .p0_rd_en   (_T_471),	// matmul/matmul-hw.mlir:20321:13
    .p1_wr_en   (_T_475),	// matmul/matmul-hw.mlir:20308:13
    .p1_wr_data (_T_474),	// matmul/matmul-hw.mlir:20309:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2274)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3632 (	// matmul/matmul-hw.mlir:20039:37
    .p0_rd_en   (_T_466),	// matmul/matmul-hw.mlir:20351:13
    .p1_wr_en   (_T_470),	// matmul/matmul-hw.mlir:20338:13
    .p1_wr_data (_T_469),	// matmul/matmul-hw.mlir:20339:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2273)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3633 (	// matmul/matmul-hw.mlir:20040:37
    .p0_rd_en   (_T_461),	// matmul/matmul-hw.mlir:20381:13
    .p1_wr_en   (_T_465),	// matmul/matmul-hw.mlir:20368:13
    .p1_wr_data (_T_464),	// matmul/matmul-hw.mlir:20369:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2272)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3634 (	// matmul/matmul-hw.mlir:20041:37
    .p0_rd_en   (_T_456),	// matmul/matmul-hw.mlir:20411:13
    .p1_wr_en   (_T_460),	// matmul/matmul-hw.mlir:20398:13
    .p1_wr_data (_T_459),	// matmul/matmul-hw.mlir:20399:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2271)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3635 (	// matmul/matmul-hw.mlir:20042:37
    .p0_rd_en   (_T_451),	// matmul/matmul-hw.mlir:20441:13
    .p1_wr_en   (_T_455),	// matmul/matmul-hw.mlir:20428:13
    .p1_wr_data (_T_454),	// matmul/matmul-hw.mlir:20429:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2270)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3636 (	// matmul/matmul-hw.mlir:20043:37
    .p0_rd_en   (_T_446),	// matmul/matmul-hw.mlir:20471:13
    .p1_wr_en   (_T_450),	// matmul/matmul-hw.mlir:20458:13
    .p1_wr_data (_T_449),	// matmul/matmul-hw.mlir:20459:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2269)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3637 (	// matmul/matmul-hw.mlir:20044:37
    .p0_rd_en   (_T_441),	// matmul/matmul-hw.mlir:20501:13
    .p1_wr_en   (_T_445),	// matmul/matmul-hw.mlir:20488:13
    .p1_wr_data (_T_444),	// matmul/matmul-hw.mlir:20489:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2268)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3638 (	// matmul/matmul-hw.mlir:20045:37
    .p0_rd_en   (_T_438),	// matmul/matmul-hw.mlir:20528:13
    .p1_wr_en   (_T_440),	// matmul/matmul-hw.mlir:20518:13
    .p1_wr_data (_T_439),	// matmul/matmul-hw.mlir:20519:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2267)
  );
  assign _T_520 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20046:13
  assign _T_519 = _T_2852 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8554:18, :20047:13
  assign _T_518 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20048:13
  assign _T_517 = _T_2841 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20049:13
  mult mult_inst160 (	// matmul/matmul-hw.mlir:20050:28
    .a      (A_reg_bank160_p0_rd_data),	// matmul/matmul-hw.mlir:12375:33
    .b      (_T_2464),
    .t      (_T_2841),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst160_result)
  );
  assign _T_516 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20051:13
  assign a_i_k_0_i_j_10 = A_reg_bank160_p0_rd_data;	// matmul/matmul-hw.mlir:12375:33, :20053:5
  //PROBE: a_i_k_0_i_j_10	// matmul/matmul-hw.mlir:20054:5
  assign b_i_k_0_i_j_10 = _T_2464;	// matmul/matmul-hw.mlir:20056:5
  //PROBE: b_i_k_0_i_j_10	// matmul/matmul-hw.mlir:20057:5
  assign c_prev_i_k_0_i_j_10 = C_reg_bank0_p0_rd_data_2283;	// matmul/matmul-hw.mlir:20029:36, :20059:5
  //PROBE: c_prev_i_k_0_i_j_10	// matmul/matmul-hw.mlir:20060:5
  assign tk_i_k_0_i_j_10 = _T_2819;	// matmul/matmul-hw.mlir:20062:5
  //PROBE: tk_i_k_0_i_j_10	// matmul/matmul-hw.mlir:20063:5
  wire [31:0] _T_3639 = mult_inst160_result + C_reg_bank0_p0_rd_data_2283;	// matmul/matmul-hw.mlir:20029:36, :20050:28, :20064:13
  assign c_i_k_0_i_j_10 = _T_3639;	// matmul/matmul-hw.mlir:20066:5
  //PROBE: c_i_k_0_i_j_10	// matmul/matmul-hw.mlir:20067:5
  assign _T_515 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20068:13
  assign _T_514 = _T_2863 ? _T_3639 : 32'bx;	// matmul/matmul-hw.mlir:8549:18, :20069:13
  localparam [3:0] _T_3641 = 4'h0;	// matmul/matmul-hw.mlir:20072:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20073:5
    if (rst)	// matmul/matmul-hw.mlir:20073:5
      i_k_next_3640 <= _T_3641;	// matmul/matmul-hw.mlir:20076:7
    else	// matmul/matmul-hw.mlir:20073:5
      i_k_next_3640 <= i_j_next_3620;	// matmul/matmul-hw.mlir:19954:13, :20074:7
  end // always @(posedge)
  assign _T_513 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20078:13
  assign _T_512 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20079:13
  mult mult_inst161 (	// matmul/matmul-hw.mlir:20080:28
    .a      (A_reg_bank161_p0_rd_data),	// matmul/matmul-hw.mlir:12376:33
    .b      (_T_2480),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst161_result)
  );
  assign _T_511 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20081:13
  assign a_i_k_1_i_j_10 = A_reg_bank161_p0_rd_data;	// matmul/matmul-hw.mlir:12376:33, :20083:5
  //PROBE: a_i_k_1_i_j_10	// matmul/matmul-hw.mlir:20084:5
  assign b_i_k_1_i_j_10 = _T_2480;	// matmul/matmul-hw.mlir:20086:5
  //PROBE: b_i_k_1_i_j_10	// matmul/matmul-hw.mlir:20087:5
  assign c_prev_i_k_1_i_j_10 = C_reg_bank1_p0_rd_data_2282;	// matmul/matmul-hw.mlir:20030:36, :20089:5
  //PROBE: c_prev_i_k_1_i_j_10	// matmul/matmul-hw.mlir:20090:5
  assign tk_i_k_1_i_j_10 = _T_2830;	// matmul/matmul-hw.mlir:20092:5
  //PROBE: tk_i_k_1_i_j_10	// matmul/matmul-hw.mlir:20093:5
  wire [31:0] _T_3642 = mult_inst161_result + C_reg_bank1_p0_rd_data_2282;	// matmul/matmul-hw.mlir:20030:36, :20080:28, :20094:13
  assign c_i_k_1_i_j_10 = _T_3642;	// matmul/matmul-hw.mlir:20096:5
  //PROBE: c_i_k_1_i_j_10	// matmul/matmul-hw.mlir:20097:5
  assign _T_510 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20098:13
  assign _T_509 = _T_2874 ? _T_3642 : 32'bx;	// matmul/matmul-hw.mlir:8544:18, :20099:13
  localparam [3:0] _T_3644 = 4'h0;	// matmul/matmul-hw.mlir:20102:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20103:5
    if (rst)	// matmul/matmul-hw.mlir:20103:5
      i_k_next_3643 <= _T_3644;	// matmul/matmul-hw.mlir:20106:7
    else	// matmul/matmul-hw.mlir:20103:5
      i_k_next_3643 <= i_k_next_3640;	// matmul/matmul-hw.mlir:20071:13, :20104:7
  end // always @(posedge)
  assign _T_508 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20108:13
  assign _T_507 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20109:13
  mult mult_inst162 (	// matmul/matmul-hw.mlir:20110:28
    .a      (A_reg_bank162_p0_rd_data),	// matmul/matmul-hw.mlir:12377:33
    .b      (_T_2496),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst162_result)
  );
  assign _T_506 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20111:13
  assign a_i_k_2_i_j_10 = A_reg_bank162_p0_rd_data;	// matmul/matmul-hw.mlir:12377:33, :20113:5
  //PROBE: a_i_k_2_i_j_10	// matmul/matmul-hw.mlir:20114:5
  assign b_i_k_2_i_j_10 = _T_2496;	// matmul/matmul-hw.mlir:20116:5
  //PROBE: b_i_k_2_i_j_10	// matmul/matmul-hw.mlir:20117:5
  assign c_prev_i_k_2_i_j_10 = C_reg_bank2_p0_rd_data_2281;	// matmul/matmul-hw.mlir:20031:36, :20119:5
  //PROBE: c_prev_i_k_2_i_j_10	// matmul/matmul-hw.mlir:20120:5
  assign tk_i_k_2_i_j_10 = _T_2841;	// matmul/matmul-hw.mlir:20122:5
  //PROBE: tk_i_k_2_i_j_10	// matmul/matmul-hw.mlir:20123:5
  wire [31:0] _T_3645 = mult_inst162_result + C_reg_bank2_p0_rd_data_2281;	// matmul/matmul-hw.mlir:20031:36, :20110:28, :20124:13
  assign c_i_k_2_i_j_10 = _T_3645;	// matmul/matmul-hw.mlir:20126:5
  //PROBE: c_i_k_2_i_j_10	// matmul/matmul-hw.mlir:20127:5
  assign _T_505 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20128:13
  assign _T_504 = _T_2885 ? _T_3645 : 32'bx;	// matmul/matmul-hw.mlir:8539:18, :20129:13
  localparam [3:0] _T_3647 = 4'h0;	// matmul/matmul-hw.mlir:20132:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20133:5
    if (rst)	// matmul/matmul-hw.mlir:20133:5
      i_k_next_3646 <= _T_3647;	// matmul/matmul-hw.mlir:20136:7
    else	// matmul/matmul-hw.mlir:20133:5
      i_k_next_3646 <= i_k_next_3643;	// matmul/matmul-hw.mlir:20101:13, :20134:7
  end // always @(posedge)
  assign _T_503 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20138:13
  assign _T_502 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20139:13
  mult mult_inst163 (	// matmul/matmul-hw.mlir:20140:28
    .a      (A_reg_bank163_p0_rd_data),	// matmul/matmul-hw.mlir:12378:33
    .b      (_T_2512),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst163_result)
  );
  assign _T_501 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20141:13
  assign a_i_k_3_i_j_10 = A_reg_bank163_p0_rd_data;	// matmul/matmul-hw.mlir:12378:33, :20143:5
  //PROBE: a_i_k_3_i_j_10	// matmul/matmul-hw.mlir:20144:5
  assign b_i_k_3_i_j_10 = _T_2512;	// matmul/matmul-hw.mlir:20146:5
  //PROBE: b_i_k_3_i_j_10	// matmul/matmul-hw.mlir:20147:5
  assign c_prev_i_k_3_i_j_10 = C_reg_bank3_p0_rd_data_2280;	// matmul/matmul-hw.mlir:20032:36, :20149:5
  //PROBE: c_prev_i_k_3_i_j_10	// matmul/matmul-hw.mlir:20150:5
  assign tk_i_k_3_i_j_10 = _T_2852;	// matmul/matmul-hw.mlir:20152:5
  //PROBE: tk_i_k_3_i_j_10	// matmul/matmul-hw.mlir:20153:5
  wire [31:0] _T_3648 = mult_inst163_result + C_reg_bank3_p0_rd_data_2280;	// matmul/matmul-hw.mlir:20032:36, :20140:28, :20154:13
  assign c_i_k_3_i_j_10 = _T_3648;	// matmul/matmul-hw.mlir:20156:5
  //PROBE: c_i_k_3_i_j_10	// matmul/matmul-hw.mlir:20157:5
  assign _T_500 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20158:13
  assign _T_499 = _T_2892 ? _T_3648 : 32'bx;	// matmul/matmul-hw.mlir:8534:18, :20159:13
  localparam [3:0] _T_3650 = 4'h0;	// matmul/matmul-hw.mlir:20162:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20163:5
    if (rst)	// matmul/matmul-hw.mlir:20163:5
      i_k_next_3649 <= _T_3650;	// matmul/matmul-hw.mlir:20166:7
    else	// matmul/matmul-hw.mlir:20163:5
      i_k_next_3649 <= i_k_next_3646;	// matmul/matmul-hw.mlir:20131:13, :20164:7
  end // always @(posedge)
  assign _T_498 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20168:13
  assign _T_497 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20169:13
  mult mult_inst164 (	// matmul/matmul-hw.mlir:20170:28
    .a      (A_reg_bank164_p0_rd_data),	// matmul/matmul-hw.mlir:12379:33
    .b      (_T_2528),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst164_result)
  );
  assign _T_496 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20171:13
  assign a_i_k_4_i_j_10 = A_reg_bank164_p0_rd_data;	// matmul/matmul-hw.mlir:12379:33, :20173:5
  //PROBE: a_i_k_4_i_j_10	// matmul/matmul-hw.mlir:20174:5
  assign b_i_k_4_i_j_10 = _T_2528;	// matmul/matmul-hw.mlir:20176:5
  //PROBE: b_i_k_4_i_j_10	// matmul/matmul-hw.mlir:20177:5
  assign c_prev_i_k_4_i_j_10 = C_reg_bank4_p0_rd_data_2279;	// matmul/matmul-hw.mlir:20033:36, :20179:5
  //PROBE: c_prev_i_k_4_i_j_10	// matmul/matmul-hw.mlir:20180:5
  assign tk_i_k_4_i_j_10 = _T_2863;	// matmul/matmul-hw.mlir:20182:5
  //PROBE: tk_i_k_4_i_j_10	// matmul/matmul-hw.mlir:20183:5
  wire [31:0] _T_3651 = mult_inst164_result + C_reg_bank4_p0_rd_data_2279;	// matmul/matmul-hw.mlir:20033:36, :20170:28, :20184:13
  assign c_i_k_4_i_j_10 = _T_3651;	// matmul/matmul-hw.mlir:20186:5
  //PROBE: c_i_k_4_i_j_10	// matmul/matmul-hw.mlir:20187:5
  assign _T_495 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20188:13
  assign _T_494 = _T_2897 ? _T_3651 : 32'bx;	// matmul/matmul-hw.mlir:8529:18, :20189:13
  localparam [3:0] _T_3653 = 4'h0;	// matmul/matmul-hw.mlir:20192:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20193:5
    if (rst)	// matmul/matmul-hw.mlir:20193:5
      i_k_next_3652 <= _T_3653;	// matmul/matmul-hw.mlir:20196:7
    else	// matmul/matmul-hw.mlir:20193:5
      i_k_next_3652 <= i_k_next_3649;	// matmul/matmul-hw.mlir:20161:13, :20194:7
  end // always @(posedge)
  assign _T_493 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20198:13
  assign _T_492 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20199:13
  mult mult_inst165 (	// matmul/matmul-hw.mlir:20200:28
    .a      (A_reg_bank165_p0_rd_data),	// matmul/matmul-hw.mlir:12380:33
    .b      (_T_2544),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst165_result)
  );
  assign _T_491 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20201:13
  assign a_i_k_5_i_j_10 = A_reg_bank165_p0_rd_data;	// matmul/matmul-hw.mlir:12380:33, :20203:5
  //PROBE: a_i_k_5_i_j_10	// matmul/matmul-hw.mlir:20204:5
  assign b_i_k_5_i_j_10 = _T_2544;	// matmul/matmul-hw.mlir:20206:5
  //PROBE: b_i_k_5_i_j_10	// matmul/matmul-hw.mlir:20207:5
  assign c_prev_i_k_5_i_j_10 = C_reg_bank5_p0_rd_data_2278;	// matmul/matmul-hw.mlir:20034:36, :20209:5
  //PROBE: c_prev_i_k_5_i_j_10	// matmul/matmul-hw.mlir:20210:5
  assign tk_i_k_5_i_j_10 = _T_2874;	// matmul/matmul-hw.mlir:20212:5
  //PROBE: tk_i_k_5_i_j_10	// matmul/matmul-hw.mlir:20213:5
  wire [31:0] _T_3654 = mult_inst165_result + C_reg_bank5_p0_rd_data_2278;	// matmul/matmul-hw.mlir:20034:36, :20200:28, :20214:13
  assign c_i_k_5_i_j_10 = _T_3654;	// matmul/matmul-hw.mlir:20216:5
  //PROBE: c_i_k_5_i_j_10	// matmul/matmul-hw.mlir:20217:5
  assign _T_490 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20218:13
  assign _T_489 = _T_2902 ? _T_3654 : 32'bx;	// matmul/matmul-hw.mlir:8524:18, :20219:13
  localparam [3:0] _T_3656 = 4'h0;	// matmul/matmul-hw.mlir:20222:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20223:5
    if (rst)	// matmul/matmul-hw.mlir:20223:5
      i_k_next_3655 <= _T_3656;	// matmul/matmul-hw.mlir:20226:7
    else	// matmul/matmul-hw.mlir:20223:5
      i_k_next_3655 <= i_k_next_3652;	// matmul/matmul-hw.mlir:20191:13, :20224:7
  end // always @(posedge)
  assign _T_488 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20228:13
  assign _T_487 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20229:13
  mult mult_inst166 (	// matmul/matmul-hw.mlir:20230:28
    .a      (A_reg_bank166_p0_rd_data),	// matmul/matmul-hw.mlir:12381:33
    .b      (_T_2560),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst166_result)
  );
  assign _T_486 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20231:13
  assign a_i_k_6_i_j_10 = A_reg_bank166_p0_rd_data;	// matmul/matmul-hw.mlir:12381:33, :20233:5
  //PROBE: a_i_k_6_i_j_10	// matmul/matmul-hw.mlir:20234:5
  assign b_i_k_6_i_j_10 = _T_2560;	// matmul/matmul-hw.mlir:20236:5
  //PROBE: b_i_k_6_i_j_10	// matmul/matmul-hw.mlir:20237:5
  assign c_prev_i_k_6_i_j_10 = C_reg_bank6_p0_rd_data_2277;	// matmul/matmul-hw.mlir:20035:36, :20239:5
  //PROBE: c_prev_i_k_6_i_j_10	// matmul/matmul-hw.mlir:20240:5
  assign tk_i_k_6_i_j_10 = _T_2885;	// matmul/matmul-hw.mlir:20242:5
  //PROBE: tk_i_k_6_i_j_10	// matmul/matmul-hw.mlir:20243:5
  wire [31:0] _T_3657 = mult_inst166_result + C_reg_bank6_p0_rd_data_2277;	// matmul/matmul-hw.mlir:20035:36, :20230:28, :20244:13
  assign c_i_k_6_i_j_10 = _T_3657;	// matmul/matmul-hw.mlir:20246:5
  //PROBE: c_i_k_6_i_j_10	// matmul/matmul-hw.mlir:20247:5
  assign _T_485 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20248:13
  assign _T_484 = _T_2907 ? _T_3657 : 32'bx;	// matmul/matmul-hw.mlir:8519:18, :20249:13
  localparam [3:0] _T_3659 = 4'h0;	// matmul/matmul-hw.mlir:20252:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20253:5
    if (rst)	// matmul/matmul-hw.mlir:20253:5
      i_k_next_3658 <= _T_3659;	// matmul/matmul-hw.mlir:20256:7
    else	// matmul/matmul-hw.mlir:20253:5
      i_k_next_3658 <= i_k_next_3655;	// matmul/matmul-hw.mlir:20221:13, :20254:7
  end // always @(posedge)
  assign _T_483 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20258:13
  assign _T_482 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20259:13
  mult mult_inst167 (	// matmul/matmul-hw.mlir:20260:28
    .a      (A_reg_bank167_p0_rd_data),	// matmul/matmul-hw.mlir:12382:33
    .b      (_T_2576),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst167_result)
  );
  assign _T_481 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20261:13
  assign a_i_k_7_i_j_10 = A_reg_bank167_p0_rd_data;	// matmul/matmul-hw.mlir:12382:33, :20263:5
  //PROBE: a_i_k_7_i_j_10	// matmul/matmul-hw.mlir:20264:5
  assign b_i_k_7_i_j_10 = _T_2576;	// matmul/matmul-hw.mlir:20266:5
  //PROBE: b_i_k_7_i_j_10	// matmul/matmul-hw.mlir:20267:5
  assign c_prev_i_k_7_i_j_10 = C_reg_bank7_p0_rd_data_2276;	// matmul/matmul-hw.mlir:20036:36, :20269:5
  //PROBE: c_prev_i_k_7_i_j_10	// matmul/matmul-hw.mlir:20270:5
  assign tk_i_k_7_i_j_10 = _T_2892;	// matmul/matmul-hw.mlir:20272:5
  //PROBE: tk_i_k_7_i_j_10	// matmul/matmul-hw.mlir:20273:5
  wire [31:0] _T_3660 = mult_inst167_result + C_reg_bank7_p0_rd_data_2276;	// matmul/matmul-hw.mlir:20036:36, :20260:28, :20274:13
  assign c_i_k_7_i_j_10 = _T_3660;	// matmul/matmul-hw.mlir:20276:5
  //PROBE: c_i_k_7_i_j_10	// matmul/matmul-hw.mlir:20277:5
  assign _T_480 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20278:13
  assign _T_479 = _T_2912 ? _T_3660 : 32'bx;	// matmul/matmul-hw.mlir:8514:18, :20279:13
  localparam [3:0] _T_3662 = 4'h0;	// matmul/matmul-hw.mlir:20282:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20283:5
    if (rst)	// matmul/matmul-hw.mlir:20283:5
      i_k_next_3661 <= _T_3662;	// matmul/matmul-hw.mlir:20286:7
    else	// matmul/matmul-hw.mlir:20283:5
      i_k_next_3661 <= i_k_next_3658;	// matmul/matmul-hw.mlir:20251:13, :20284:7
  end // always @(posedge)
  assign _T_478 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20288:13
  assign _T_477 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20289:13
  mult mult_inst168 (	// matmul/matmul-hw.mlir:20290:28
    .a      (A_reg_bank168_p0_rd_data),	// matmul/matmul-hw.mlir:12383:33
    .b      (_T_2592),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst168_result)
  );
  assign _T_476 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20291:13
  assign a_i_k_8_i_j_10 = A_reg_bank168_p0_rd_data;	// matmul/matmul-hw.mlir:12383:33, :20293:5
  //PROBE: a_i_k_8_i_j_10	// matmul/matmul-hw.mlir:20294:5
  assign b_i_k_8_i_j_10 = _T_2592;	// matmul/matmul-hw.mlir:20296:5
  //PROBE: b_i_k_8_i_j_10	// matmul/matmul-hw.mlir:20297:5
  assign c_prev_i_k_8_i_j_10 = C_reg_bank8_p0_rd_data_2275;	// matmul/matmul-hw.mlir:20037:36, :20299:5
  //PROBE: c_prev_i_k_8_i_j_10	// matmul/matmul-hw.mlir:20300:5
  assign tk_i_k_8_i_j_10 = _T_2897;	// matmul/matmul-hw.mlir:20302:5
  //PROBE: tk_i_k_8_i_j_10	// matmul/matmul-hw.mlir:20303:5
  wire [31:0] _T_3663 = mult_inst168_result + C_reg_bank8_p0_rd_data_2275;	// matmul/matmul-hw.mlir:20037:36, :20290:28, :20304:13
  assign c_i_k_8_i_j_10 = _T_3663;	// matmul/matmul-hw.mlir:20306:5
  //PROBE: c_i_k_8_i_j_10	// matmul/matmul-hw.mlir:20307:5
  assign _T_475 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20308:13
  assign _T_474 = _T_2917 ? _T_3663 : 32'bx;	// matmul/matmul-hw.mlir:8509:18, :20309:13
  localparam [3:0] _T_3665 = 4'h0;	// matmul/matmul-hw.mlir:20312:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20313:5
    if (rst)	// matmul/matmul-hw.mlir:20313:5
      i_k_next_3664 <= _T_3665;	// matmul/matmul-hw.mlir:20316:7
    else	// matmul/matmul-hw.mlir:20313:5
      i_k_next_3664 <= i_k_next_3661;	// matmul/matmul-hw.mlir:20281:13, :20314:7
  end // always @(posedge)
  assign _T_473 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20318:13
  assign _T_472 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20319:13
  mult mult_inst169 (	// matmul/matmul-hw.mlir:20320:28
    .a      (A_reg_bank169_p0_rd_data),	// matmul/matmul-hw.mlir:12384:33
    .b      (_T_2608),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst169_result)
  );
  assign _T_471 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20321:13
  assign a_i_k_9_i_j_10 = A_reg_bank169_p0_rd_data;	// matmul/matmul-hw.mlir:12384:33, :20323:5
  //PROBE: a_i_k_9_i_j_10	// matmul/matmul-hw.mlir:20324:5
  assign b_i_k_9_i_j_10 = _T_2608;	// matmul/matmul-hw.mlir:20326:5
  //PROBE: b_i_k_9_i_j_10	// matmul/matmul-hw.mlir:20327:5
  assign c_prev_i_k_9_i_j_10 = C_reg_bank9_p0_rd_data_2274;	// matmul/matmul-hw.mlir:20038:36, :20329:5
  //PROBE: c_prev_i_k_9_i_j_10	// matmul/matmul-hw.mlir:20330:5
  assign tk_i_k_9_i_j_10 = _T_2902;	// matmul/matmul-hw.mlir:20332:5
  //PROBE: tk_i_k_9_i_j_10	// matmul/matmul-hw.mlir:20333:5
  wire [31:0] _T_3666 = mult_inst169_result + C_reg_bank9_p0_rd_data_2274;	// matmul/matmul-hw.mlir:20038:36, :20320:28, :20334:13
  assign c_i_k_9_i_j_10 = _T_3666;	// matmul/matmul-hw.mlir:20336:5
  //PROBE: c_i_k_9_i_j_10	// matmul/matmul-hw.mlir:20337:5
  assign _T_470 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20338:13
  assign _T_469 = _T_2922 ? _T_3666 : 32'bx;	// matmul/matmul-hw.mlir:8504:18, :20339:13
  localparam [3:0] _T_3668 = 4'h0;	// matmul/matmul-hw.mlir:20342:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20343:5
    if (rst)	// matmul/matmul-hw.mlir:20343:5
      i_k_next_3667 <= _T_3668;	// matmul/matmul-hw.mlir:20346:7
    else	// matmul/matmul-hw.mlir:20343:5
      i_k_next_3667 <= i_k_next_3664;	// matmul/matmul-hw.mlir:20311:13, :20344:7
  end // always @(posedge)
  assign _T_468 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20348:13
  assign _T_467 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20349:13
  mult mult_inst170 (	// matmul/matmul-hw.mlir:20350:28
    .a      (A_reg_bank170_p0_rd_data),	// matmul/matmul-hw.mlir:12385:33
    .b      (_T_2624),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst170_result)
  );
  assign _T_466 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20351:13
  assign a_i_k_10_i_j_10 = A_reg_bank170_p0_rd_data;	// matmul/matmul-hw.mlir:12385:33, :20353:5
  //PROBE: a_i_k_10_i_j_10	// matmul/matmul-hw.mlir:20354:5
  assign b_i_k_10_i_j_10 = _T_2624;	// matmul/matmul-hw.mlir:20356:5
  //PROBE: b_i_k_10_i_j_10	// matmul/matmul-hw.mlir:20357:5
  assign c_prev_i_k_10_i_j_10 = C_reg_bank10_p0_rd_data_2273;	// matmul/matmul-hw.mlir:20039:37, :20359:5
  //PROBE: c_prev_i_k_10_i_j_10	// matmul/matmul-hw.mlir:20360:5
  assign tk_i_k_10_i_j_10 = _T_2907;	// matmul/matmul-hw.mlir:20362:5
  //PROBE: tk_i_k_10_i_j_10	// matmul/matmul-hw.mlir:20363:5
  wire [31:0] _T_3669 = mult_inst170_result + C_reg_bank10_p0_rd_data_2273;	// matmul/matmul-hw.mlir:20039:37, :20350:28, :20364:13
  assign c_i_k_10_i_j_10 = _T_3669;	// matmul/matmul-hw.mlir:20366:5
  //PROBE: c_i_k_10_i_j_10	// matmul/matmul-hw.mlir:20367:5
  assign _T_465 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20368:13
  assign _T_464 = _T_2927 ? _T_3669 : 32'bx;	// matmul/matmul-hw.mlir:8499:18, :20369:13
  localparam [3:0] _T_3671 = 4'h0;	// matmul/matmul-hw.mlir:20372:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20373:5
    if (rst)	// matmul/matmul-hw.mlir:20373:5
      i_k_next_3670 <= _T_3671;	// matmul/matmul-hw.mlir:20376:7
    else	// matmul/matmul-hw.mlir:20373:5
      i_k_next_3670 <= i_k_next_3667;	// matmul/matmul-hw.mlir:20341:13, :20374:7
  end // always @(posedge)
  assign _T_463 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20378:13
  assign _T_462 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20379:13
  mult mult_inst171 (	// matmul/matmul-hw.mlir:20380:28
    .a      (A_reg_bank171_p0_rd_data),	// matmul/matmul-hw.mlir:12386:33
    .b      (_T_2640),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst171_result)
  );
  assign _T_461 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20381:13
  assign a_i_k_11_i_j_10 = A_reg_bank171_p0_rd_data;	// matmul/matmul-hw.mlir:12386:33, :20383:5
  //PROBE: a_i_k_11_i_j_10	// matmul/matmul-hw.mlir:20384:5
  assign b_i_k_11_i_j_10 = _T_2640;	// matmul/matmul-hw.mlir:20386:5
  //PROBE: b_i_k_11_i_j_10	// matmul/matmul-hw.mlir:20387:5
  assign c_prev_i_k_11_i_j_10 = C_reg_bank11_p0_rd_data_2272;	// matmul/matmul-hw.mlir:20040:37, :20389:5
  //PROBE: c_prev_i_k_11_i_j_10	// matmul/matmul-hw.mlir:20390:5
  assign tk_i_k_11_i_j_10 = _T_2912;	// matmul/matmul-hw.mlir:20392:5
  //PROBE: tk_i_k_11_i_j_10	// matmul/matmul-hw.mlir:20393:5
  wire [31:0] _T_3672 = mult_inst171_result + C_reg_bank11_p0_rd_data_2272;	// matmul/matmul-hw.mlir:20040:37, :20380:28, :20394:13
  assign c_i_k_11_i_j_10 = _T_3672;	// matmul/matmul-hw.mlir:20396:5
  //PROBE: c_i_k_11_i_j_10	// matmul/matmul-hw.mlir:20397:5
  assign _T_460 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20398:13
  assign _T_459 = _T_2932 ? _T_3672 : 32'bx;	// matmul/matmul-hw.mlir:8494:18, :20399:13
  localparam [3:0] _T_3674 = 4'h0;	// matmul/matmul-hw.mlir:20402:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20403:5
    if (rst)	// matmul/matmul-hw.mlir:20403:5
      i_k_next_3673 <= _T_3674;	// matmul/matmul-hw.mlir:20406:7
    else	// matmul/matmul-hw.mlir:20403:5
      i_k_next_3673 <= i_k_next_3670;	// matmul/matmul-hw.mlir:20371:13, :20404:7
  end // always @(posedge)
  assign _T_458 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20408:13
  assign _T_457 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20409:13
  mult mult_inst172 (	// matmul/matmul-hw.mlir:20410:28
    .a      (A_reg_bank172_p0_rd_data),	// matmul/matmul-hw.mlir:12387:33
    .b      (_T_2656),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst172_result)
  );
  assign _T_456 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20411:13
  assign a_i_k_12_i_j_10 = A_reg_bank172_p0_rd_data;	// matmul/matmul-hw.mlir:12387:33, :20413:5
  //PROBE: a_i_k_12_i_j_10	// matmul/matmul-hw.mlir:20414:5
  assign b_i_k_12_i_j_10 = _T_2656;	// matmul/matmul-hw.mlir:20416:5
  //PROBE: b_i_k_12_i_j_10	// matmul/matmul-hw.mlir:20417:5
  assign c_prev_i_k_12_i_j_10 = C_reg_bank12_p0_rd_data_2271;	// matmul/matmul-hw.mlir:20041:37, :20419:5
  //PROBE: c_prev_i_k_12_i_j_10	// matmul/matmul-hw.mlir:20420:5
  assign tk_i_k_12_i_j_10 = _T_2917;	// matmul/matmul-hw.mlir:20422:5
  //PROBE: tk_i_k_12_i_j_10	// matmul/matmul-hw.mlir:20423:5
  wire [31:0] _T_3675 = mult_inst172_result + C_reg_bank12_p0_rd_data_2271;	// matmul/matmul-hw.mlir:20041:37, :20410:28, :20424:13
  assign c_i_k_12_i_j_10 = _T_3675;	// matmul/matmul-hw.mlir:20426:5
  //PROBE: c_i_k_12_i_j_10	// matmul/matmul-hw.mlir:20427:5
  assign _T_455 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20428:13
  assign _T_454 = _T_2937 ? _T_3675 : 32'bx;	// matmul/matmul-hw.mlir:8489:18, :20429:13
  localparam [3:0] _T_3677 = 4'h0;	// matmul/matmul-hw.mlir:20432:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20433:5
    if (rst)	// matmul/matmul-hw.mlir:20433:5
      i_k_next_3676 <= _T_3677;	// matmul/matmul-hw.mlir:20436:7
    else	// matmul/matmul-hw.mlir:20433:5
      i_k_next_3676 <= i_k_next_3673;	// matmul/matmul-hw.mlir:20401:13, :20434:7
  end // always @(posedge)
  assign _T_453 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20438:13
  assign _T_452 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20439:13
  mult mult_inst173 (	// matmul/matmul-hw.mlir:20440:28
    .a      (A_reg_bank173_p0_rd_data),	// matmul/matmul-hw.mlir:12388:33
    .b      (_T_2672),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst173_result)
  );
  assign _T_451 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20441:13
  assign a_i_k_13_i_j_10 = A_reg_bank173_p0_rd_data;	// matmul/matmul-hw.mlir:12388:33, :20443:5
  //PROBE: a_i_k_13_i_j_10	// matmul/matmul-hw.mlir:20444:5
  assign b_i_k_13_i_j_10 = _T_2672;	// matmul/matmul-hw.mlir:20446:5
  //PROBE: b_i_k_13_i_j_10	// matmul/matmul-hw.mlir:20447:5
  assign c_prev_i_k_13_i_j_10 = C_reg_bank13_p0_rd_data_2270;	// matmul/matmul-hw.mlir:20042:37, :20449:5
  //PROBE: c_prev_i_k_13_i_j_10	// matmul/matmul-hw.mlir:20450:5
  assign tk_i_k_13_i_j_10 = _T_2922;	// matmul/matmul-hw.mlir:20452:5
  //PROBE: tk_i_k_13_i_j_10	// matmul/matmul-hw.mlir:20453:5
  wire [31:0] _T_3678 = mult_inst173_result + C_reg_bank13_p0_rd_data_2270;	// matmul/matmul-hw.mlir:20042:37, :20440:28, :20454:13
  assign c_i_k_13_i_j_10 = _T_3678;	// matmul/matmul-hw.mlir:20456:5
  //PROBE: c_i_k_13_i_j_10	// matmul/matmul-hw.mlir:20457:5
  assign _T_450 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20458:13
  assign _T_449 = _T_2942 ? _T_3678 : 32'bx;	// matmul/matmul-hw.mlir:8484:18, :20459:13
  localparam [3:0] _T_3680 = 4'h0;	// matmul/matmul-hw.mlir:20462:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20463:5
    if (rst)	// matmul/matmul-hw.mlir:20463:5
      i_k_next_3679 <= _T_3680;	// matmul/matmul-hw.mlir:20466:7
    else	// matmul/matmul-hw.mlir:20463:5
      i_k_next_3679 <= i_k_next_3676;	// matmul/matmul-hw.mlir:20431:13, :20464:7
  end // always @(posedge)
  assign _T_448 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20468:13
  assign _T_447 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20469:13
  mult mult_inst174 (	// matmul/matmul-hw.mlir:20470:28
    .a      (A_reg_bank174_p0_rd_data),	// matmul/matmul-hw.mlir:12389:33
    .b      (_T_2688),
    .t      (_T_2937),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst174_result)
  );
  assign _T_446 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20471:13
  assign a_i_k_14_i_j_10 = A_reg_bank174_p0_rd_data;	// matmul/matmul-hw.mlir:12389:33, :20473:5
  //PROBE: a_i_k_14_i_j_10	// matmul/matmul-hw.mlir:20474:5
  assign b_i_k_14_i_j_10 = _T_2688;	// matmul/matmul-hw.mlir:20476:5
  //PROBE: b_i_k_14_i_j_10	// matmul/matmul-hw.mlir:20477:5
  assign c_prev_i_k_14_i_j_10 = C_reg_bank14_p0_rd_data_2269;	// matmul/matmul-hw.mlir:20043:37, :20479:5
  //PROBE: c_prev_i_k_14_i_j_10	// matmul/matmul-hw.mlir:20480:5
  assign tk_i_k_14_i_j_10 = _T_2927;	// matmul/matmul-hw.mlir:20482:5
  //PROBE: tk_i_k_14_i_j_10	// matmul/matmul-hw.mlir:20483:5
  wire [31:0] _T_3681 = mult_inst174_result + C_reg_bank14_p0_rd_data_2269;	// matmul/matmul-hw.mlir:20043:37, :20470:28, :20484:13
  assign c_i_k_14_i_j_10 = _T_3681;	// matmul/matmul-hw.mlir:20486:5
  //PROBE: c_i_k_14_i_j_10	// matmul/matmul-hw.mlir:20487:5
  assign _T_445 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20488:13
  assign _T_444 = _T_2947 ? _T_3681 : 32'bx;	// matmul/matmul-hw.mlir:8479:18, :20489:13
  localparam [3:0] _T_3683 = 4'h0;	// matmul/matmul-hw.mlir:20492:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20493:5
    if (rst)	// matmul/matmul-hw.mlir:20493:5
      i_k_next_3682 <= _T_3683;	// matmul/matmul-hw.mlir:20496:7
    else	// matmul/matmul-hw.mlir:20493:5
      i_k_next_3682 <= i_k_next_3679;	// matmul/matmul-hw.mlir:20461:13, :20494:7
  end // always @(posedge)
  assign _T_443 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20498:13
  assign _T_442 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20499:13
  mult mult_inst175 (	// matmul/matmul-hw.mlir:20500:28
    .a      (A_reg_bank175_p0_rd_data),	// matmul/matmul-hw.mlir:12390:33
    .b      (_T_2704),
    .t      (_T_2942),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst175_result)
  );
  assign _T_441 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20501:13
  assign a_i_k_15_i_j_10 = A_reg_bank175_p0_rd_data;	// matmul/matmul-hw.mlir:12390:33, :20503:5
  //PROBE: a_i_k_15_i_j_10	// matmul/matmul-hw.mlir:20504:5
  assign b_i_k_15_i_j_10 = _T_2704;	// matmul/matmul-hw.mlir:20506:5
  //PROBE: b_i_k_15_i_j_10	// matmul/matmul-hw.mlir:20507:5
  assign c_prev_i_k_15_i_j_10 = C_reg_bank15_p0_rd_data_2268;	// matmul/matmul-hw.mlir:20044:37, :20509:5
  //PROBE: c_prev_i_k_15_i_j_10	// matmul/matmul-hw.mlir:20510:5
  assign tk_i_k_15_i_j_10 = _T_2932;	// matmul/matmul-hw.mlir:20512:5
  //PROBE: tk_i_k_15_i_j_10	// matmul/matmul-hw.mlir:20513:5
  wire [31:0] _T_3684 = mult_inst175_result + C_reg_bank15_p0_rd_data_2268;	// matmul/matmul-hw.mlir:20044:37, :20500:28, :20514:13
  assign c_i_k_15_i_j_10 = _T_3684;	// matmul/matmul-hw.mlir:20516:5
  //PROBE: c_i_k_15_i_j_10	// matmul/matmul-hw.mlir:20517:5
  assign _T_440 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20518:13
  assign _T_439 = _T_2952 ? _T_3684 : 32'bx;	// matmul/matmul-hw.mlir:8474:18, :20519:13
  localparam [3:0] _T_3686 = 4'h0;	// matmul/matmul-hw.mlir:20522:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20523:5
    if (rst)	// matmul/matmul-hw.mlir:20523:5
      i_k_next_3685 <= _T_3686;	// matmul/matmul-hw.mlir:20526:7
    else	// matmul/matmul-hw.mlir:20523:5
      i_k_next_3685 <= i_k_next_3682;	// matmul/matmul-hw.mlir:20491:13, :20524:7
  end // always @(posedge)
  assign _T_438 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20528:13
  wire [3:0][3:0] _T_3688 = i_delayed_3687;	// matmul/matmul-hw.mlir:20530:13
  wire [3:0][3:0] _T_3689 = {_T_3688[2'h0+:3], {{i_k_next_3685}}};	// matmul/matmul-hw.mlir:20521:13, :20531:19, :20532:13, :20533:13, :20534:13
  wire [3:0][3:0] _T_3690 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:20535:19, :20536:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20537:5
    if (rst)	// matmul/matmul-hw.mlir:20537:5
      i_delayed_3687 <= _T_3690;	// matmul/matmul-hw.mlir:20540:7
    else	// matmul/matmul-hw.mlir:20537:5
      i_delayed_3687 <= _T_3689;	// matmul/matmul-hw.mlir:20538:7
  end // always @(posedge)
  assign _T_437 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20544:13
  assign _T_436 = _T_2957 ? i_delayed_3687[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8471:17, :20530:13, :20542:20, :20543:13, :20545:13
  assign _T_435 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20546:13
  assign _T_434 = _T_2957 ? C_reg_bank16_p0_rd_data_2267 : 32'bx;	// matmul/matmul-hw.mlir:8469:18, :20045:37, :20547:13
  localparam [3:0] _T_3692 = 4'h0;	// matmul/matmul-hw.mlir:20550:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20551:5
    if (rst)	// matmul/matmul-hw.mlir:20551:5
      i_j_next_3691 <= _T_3692;	// matmul/matmul-hw.mlir:20554:7
    else	// matmul/matmul-hw.mlir:20551:5
      i_j_next_3691 <= i_j_next_3620;	// matmul/matmul-hw.mlir:19954:13, :20552:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3693 (	// matmul/matmul-hw.mlir:20624:36
    .p0_rd_en   (_T_429),	// matmul/matmul-hw.mlir:20646:13
    .p1_wr_en   (_T_433),	// matmul/matmul-hw.mlir:20641:13
    .p1_wr_data (_T_432),	// matmul/matmul-hw.mlir:20642:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2266)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3694 (	// matmul/matmul-hw.mlir:20625:36
    .p0_rd_en   (_T_424),	// matmul/matmul-hw.mlir:20676:13
    .p1_wr_en   (_T_428),	// matmul/matmul-hw.mlir:20663:13
    .p1_wr_data (_T_427),	// matmul/matmul-hw.mlir:20664:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2265)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3695 (	// matmul/matmul-hw.mlir:20626:36
    .p0_rd_en   (_T_419),	// matmul/matmul-hw.mlir:20706:13
    .p1_wr_en   (_T_423),	// matmul/matmul-hw.mlir:20693:13
    .p1_wr_data (_T_422),	// matmul/matmul-hw.mlir:20694:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2264)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3696 (	// matmul/matmul-hw.mlir:20627:36
    .p0_rd_en   (_T_414),	// matmul/matmul-hw.mlir:20736:13
    .p1_wr_en   (_T_418),	// matmul/matmul-hw.mlir:20723:13
    .p1_wr_data (_T_417),	// matmul/matmul-hw.mlir:20724:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2263)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3697 (	// matmul/matmul-hw.mlir:20628:36
    .p0_rd_en   (_T_409),	// matmul/matmul-hw.mlir:20766:13
    .p1_wr_en   (_T_413),	// matmul/matmul-hw.mlir:20753:13
    .p1_wr_data (_T_412),	// matmul/matmul-hw.mlir:20754:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2262)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3698 (	// matmul/matmul-hw.mlir:20629:36
    .p0_rd_en   (_T_404),	// matmul/matmul-hw.mlir:20796:13
    .p1_wr_en   (_T_408),	// matmul/matmul-hw.mlir:20783:13
    .p1_wr_data (_T_407),	// matmul/matmul-hw.mlir:20784:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2261)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3699 (	// matmul/matmul-hw.mlir:20630:36
    .p0_rd_en   (_T_399),	// matmul/matmul-hw.mlir:20826:13
    .p1_wr_en   (_T_403),	// matmul/matmul-hw.mlir:20813:13
    .p1_wr_data (_T_402),	// matmul/matmul-hw.mlir:20814:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2260)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3700 (	// matmul/matmul-hw.mlir:20631:36
    .p0_rd_en   (_T_394),	// matmul/matmul-hw.mlir:20856:13
    .p1_wr_en   (_T_398),	// matmul/matmul-hw.mlir:20843:13
    .p1_wr_data (_T_397),	// matmul/matmul-hw.mlir:20844:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2259)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3701 (	// matmul/matmul-hw.mlir:20632:36
    .p0_rd_en   (_T_389),	// matmul/matmul-hw.mlir:20886:13
    .p1_wr_en   (_T_393),	// matmul/matmul-hw.mlir:20873:13
    .p1_wr_data (_T_392),	// matmul/matmul-hw.mlir:20874:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2258)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3702 (	// matmul/matmul-hw.mlir:20633:36
    .p0_rd_en   (_T_384),	// matmul/matmul-hw.mlir:20916:13
    .p1_wr_en   (_T_388),	// matmul/matmul-hw.mlir:20903:13
    .p1_wr_data (_T_387),	// matmul/matmul-hw.mlir:20904:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2257)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3703 (	// matmul/matmul-hw.mlir:20634:37
    .p0_rd_en   (_T_379),	// matmul/matmul-hw.mlir:20946:13
    .p1_wr_en   (_T_383),	// matmul/matmul-hw.mlir:20933:13
    .p1_wr_data (_T_382),	// matmul/matmul-hw.mlir:20934:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2256)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3704 (	// matmul/matmul-hw.mlir:20635:37
    .p0_rd_en   (_T_374),	// matmul/matmul-hw.mlir:20976:13
    .p1_wr_en   (_T_378),	// matmul/matmul-hw.mlir:20963:13
    .p1_wr_data (_T_377),	// matmul/matmul-hw.mlir:20964:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2255)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3705 (	// matmul/matmul-hw.mlir:20636:37
    .p0_rd_en   (_T_369),	// matmul/matmul-hw.mlir:21006:13
    .p1_wr_en   (_T_373),	// matmul/matmul-hw.mlir:20993:13
    .p1_wr_data (_T_372),	// matmul/matmul-hw.mlir:20994:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2254)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3706 (	// matmul/matmul-hw.mlir:20637:37
    .p0_rd_en   (_T_364),	// matmul/matmul-hw.mlir:21036:13
    .p1_wr_en   (_T_368),	// matmul/matmul-hw.mlir:21023:13
    .p1_wr_data (_T_367),	// matmul/matmul-hw.mlir:21024:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2253)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3707 (	// matmul/matmul-hw.mlir:20638:37
    .p0_rd_en   (_T_359),	// matmul/matmul-hw.mlir:21066:13
    .p1_wr_en   (_T_363),	// matmul/matmul-hw.mlir:21053:13
    .p1_wr_data (_T_362),	// matmul/matmul-hw.mlir:21054:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2252)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3708 (	// matmul/matmul-hw.mlir:20639:37
    .p0_rd_en   (_T_354),	// matmul/matmul-hw.mlir:21096:13
    .p1_wr_en   (_T_358),	// matmul/matmul-hw.mlir:21083:13
    .p1_wr_data (_T_357),	// matmul/matmul-hw.mlir:21084:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2251)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3709 (	// matmul/matmul-hw.mlir:20640:37
    .p0_rd_en   (_T_351),	// matmul/matmul-hw.mlir:21123:13
    .p1_wr_en   (_T_353),	// matmul/matmul-hw.mlir:21113:13
    .p1_wr_data (_T_352),	// matmul/matmul-hw.mlir:21114:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2250)
  );
  assign _T_433 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20641:13
  assign _T_432 = _T_2863 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8467:18, :20642:13
  assign _T_431 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20643:13
  assign _T_430 = _T_2852 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20644:13
  mult mult_inst176 (	// matmul/matmul-hw.mlir:20645:28
    .a      (A_reg_bank176_p0_rd_data),	// matmul/matmul-hw.mlir:12391:33
    .b      (_T_2465),
    .t      (_T_2852),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst176_result)
  );
  assign _T_429 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20646:13
  assign a_i_k_0_i_j_11 = A_reg_bank176_p0_rd_data;	// matmul/matmul-hw.mlir:12391:33, :20648:5
  //PROBE: a_i_k_0_i_j_11	// matmul/matmul-hw.mlir:20649:5
  assign b_i_k_0_i_j_11 = _T_2465;	// matmul/matmul-hw.mlir:20651:5
  //PROBE: b_i_k_0_i_j_11	// matmul/matmul-hw.mlir:20652:5
  assign c_prev_i_k_0_i_j_11 = C_reg_bank0_p0_rd_data_2266;	// matmul/matmul-hw.mlir:20624:36, :20654:5
  //PROBE: c_prev_i_k_0_i_j_11	// matmul/matmul-hw.mlir:20655:5
  assign tk_i_k_0_i_j_11 = _T_2830;	// matmul/matmul-hw.mlir:20657:5
  //PROBE: tk_i_k_0_i_j_11	// matmul/matmul-hw.mlir:20658:5
  wire [31:0] _T_3710 = mult_inst176_result + C_reg_bank0_p0_rd_data_2266;	// matmul/matmul-hw.mlir:20624:36, :20645:28, :20659:13
  assign c_i_k_0_i_j_11 = _T_3710;	// matmul/matmul-hw.mlir:20661:5
  //PROBE: c_i_k_0_i_j_11	// matmul/matmul-hw.mlir:20662:5
  assign _T_428 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20663:13
  assign _T_427 = _T_2874 ? _T_3710 : 32'bx;	// matmul/matmul-hw.mlir:8462:18, :20664:13
  localparam [3:0] _T_3712 = 4'h0;	// matmul/matmul-hw.mlir:20667:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20668:5
    if (rst)	// matmul/matmul-hw.mlir:20668:5
      i_k_next_3711 <= _T_3712;	// matmul/matmul-hw.mlir:20671:7
    else	// matmul/matmul-hw.mlir:20668:5
      i_k_next_3711 <= i_j_next_3691;	// matmul/matmul-hw.mlir:20549:13, :20669:7
  end // always @(posedge)
  assign _T_426 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20673:13
  assign _T_425 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20674:13
  mult mult_inst177 (	// matmul/matmul-hw.mlir:20675:28
    .a      (A_reg_bank177_p0_rd_data),	// matmul/matmul-hw.mlir:12392:33
    .b      (_T_2481),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst177_result)
  );
  assign _T_424 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20676:13
  assign a_i_k_1_i_j_11 = A_reg_bank177_p0_rd_data;	// matmul/matmul-hw.mlir:12392:33, :20678:5
  //PROBE: a_i_k_1_i_j_11	// matmul/matmul-hw.mlir:20679:5
  assign b_i_k_1_i_j_11 = _T_2481;	// matmul/matmul-hw.mlir:20681:5
  //PROBE: b_i_k_1_i_j_11	// matmul/matmul-hw.mlir:20682:5
  assign c_prev_i_k_1_i_j_11 = C_reg_bank1_p0_rd_data_2265;	// matmul/matmul-hw.mlir:20625:36, :20684:5
  //PROBE: c_prev_i_k_1_i_j_11	// matmul/matmul-hw.mlir:20685:5
  assign tk_i_k_1_i_j_11 = _T_2841;	// matmul/matmul-hw.mlir:20687:5
  //PROBE: tk_i_k_1_i_j_11	// matmul/matmul-hw.mlir:20688:5
  wire [31:0] _T_3713 = mult_inst177_result + C_reg_bank1_p0_rd_data_2265;	// matmul/matmul-hw.mlir:20625:36, :20675:28, :20689:13
  assign c_i_k_1_i_j_11 = _T_3713;	// matmul/matmul-hw.mlir:20691:5
  //PROBE: c_i_k_1_i_j_11	// matmul/matmul-hw.mlir:20692:5
  assign _T_423 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20693:13
  assign _T_422 = _T_2885 ? _T_3713 : 32'bx;	// matmul/matmul-hw.mlir:8457:18, :20694:13
  localparam [3:0] _T_3715 = 4'h0;	// matmul/matmul-hw.mlir:20697:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20698:5
    if (rst)	// matmul/matmul-hw.mlir:20698:5
      i_k_next_3714 <= _T_3715;	// matmul/matmul-hw.mlir:20701:7
    else	// matmul/matmul-hw.mlir:20698:5
      i_k_next_3714 <= i_k_next_3711;	// matmul/matmul-hw.mlir:20666:13, :20699:7
  end // always @(posedge)
  assign _T_421 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20703:13
  assign _T_420 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20704:13
  mult mult_inst178 (	// matmul/matmul-hw.mlir:20705:28
    .a      (A_reg_bank178_p0_rd_data),	// matmul/matmul-hw.mlir:12393:33
    .b      (_T_2497),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst178_result)
  );
  assign _T_419 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20706:13
  assign a_i_k_2_i_j_11 = A_reg_bank178_p0_rd_data;	// matmul/matmul-hw.mlir:12393:33, :20708:5
  //PROBE: a_i_k_2_i_j_11	// matmul/matmul-hw.mlir:20709:5
  assign b_i_k_2_i_j_11 = _T_2497;	// matmul/matmul-hw.mlir:20711:5
  //PROBE: b_i_k_2_i_j_11	// matmul/matmul-hw.mlir:20712:5
  assign c_prev_i_k_2_i_j_11 = C_reg_bank2_p0_rd_data_2264;	// matmul/matmul-hw.mlir:20626:36, :20714:5
  //PROBE: c_prev_i_k_2_i_j_11	// matmul/matmul-hw.mlir:20715:5
  assign tk_i_k_2_i_j_11 = _T_2852;	// matmul/matmul-hw.mlir:20717:5
  //PROBE: tk_i_k_2_i_j_11	// matmul/matmul-hw.mlir:20718:5
  wire [31:0] _T_3716 = mult_inst178_result + C_reg_bank2_p0_rd_data_2264;	// matmul/matmul-hw.mlir:20626:36, :20705:28, :20719:13
  assign c_i_k_2_i_j_11 = _T_3716;	// matmul/matmul-hw.mlir:20721:5
  //PROBE: c_i_k_2_i_j_11	// matmul/matmul-hw.mlir:20722:5
  assign _T_418 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20723:13
  assign _T_417 = _T_2892 ? _T_3716 : 32'bx;	// matmul/matmul-hw.mlir:8452:18, :20724:13
  localparam [3:0] _T_3718 = 4'h0;	// matmul/matmul-hw.mlir:20727:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20728:5
    if (rst)	// matmul/matmul-hw.mlir:20728:5
      i_k_next_3717 <= _T_3718;	// matmul/matmul-hw.mlir:20731:7
    else	// matmul/matmul-hw.mlir:20728:5
      i_k_next_3717 <= i_k_next_3714;	// matmul/matmul-hw.mlir:20696:13, :20729:7
  end // always @(posedge)
  assign _T_416 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20733:13
  assign _T_415 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20734:13
  mult mult_inst179 (	// matmul/matmul-hw.mlir:20735:28
    .a      (A_reg_bank179_p0_rd_data),	// matmul/matmul-hw.mlir:12394:33
    .b      (_T_2513),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst179_result)
  );
  assign _T_414 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20736:13
  assign a_i_k_3_i_j_11 = A_reg_bank179_p0_rd_data;	// matmul/matmul-hw.mlir:12394:33, :20738:5
  //PROBE: a_i_k_3_i_j_11	// matmul/matmul-hw.mlir:20739:5
  assign b_i_k_3_i_j_11 = _T_2513;	// matmul/matmul-hw.mlir:20741:5
  //PROBE: b_i_k_3_i_j_11	// matmul/matmul-hw.mlir:20742:5
  assign c_prev_i_k_3_i_j_11 = C_reg_bank3_p0_rd_data_2263;	// matmul/matmul-hw.mlir:20627:36, :20744:5
  //PROBE: c_prev_i_k_3_i_j_11	// matmul/matmul-hw.mlir:20745:5
  assign tk_i_k_3_i_j_11 = _T_2863;	// matmul/matmul-hw.mlir:20747:5
  //PROBE: tk_i_k_3_i_j_11	// matmul/matmul-hw.mlir:20748:5
  wire [31:0] _T_3719 = mult_inst179_result + C_reg_bank3_p0_rd_data_2263;	// matmul/matmul-hw.mlir:20627:36, :20735:28, :20749:13
  assign c_i_k_3_i_j_11 = _T_3719;	// matmul/matmul-hw.mlir:20751:5
  //PROBE: c_i_k_3_i_j_11	// matmul/matmul-hw.mlir:20752:5
  assign _T_413 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20753:13
  assign _T_412 = _T_2897 ? _T_3719 : 32'bx;	// matmul/matmul-hw.mlir:8447:18, :20754:13
  localparam [3:0] _T_3721 = 4'h0;	// matmul/matmul-hw.mlir:20757:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20758:5
    if (rst)	// matmul/matmul-hw.mlir:20758:5
      i_k_next_3720 <= _T_3721;	// matmul/matmul-hw.mlir:20761:7
    else	// matmul/matmul-hw.mlir:20758:5
      i_k_next_3720 <= i_k_next_3717;	// matmul/matmul-hw.mlir:20726:13, :20759:7
  end // always @(posedge)
  assign _T_411 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20763:13
  assign _T_410 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20764:13
  mult mult_inst180 (	// matmul/matmul-hw.mlir:20765:28
    .a      (A_reg_bank180_p0_rd_data),	// matmul/matmul-hw.mlir:12395:33
    .b      (_T_2529),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst180_result)
  );
  assign _T_409 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20766:13
  assign a_i_k_4_i_j_11 = A_reg_bank180_p0_rd_data;	// matmul/matmul-hw.mlir:12395:33, :20768:5
  //PROBE: a_i_k_4_i_j_11	// matmul/matmul-hw.mlir:20769:5
  assign b_i_k_4_i_j_11 = _T_2529;	// matmul/matmul-hw.mlir:20771:5
  //PROBE: b_i_k_4_i_j_11	// matmul/matmul-hw.mlir:20772:5
  assign c_prev_i_k_4_i_j_11 = C_reg_bank4_p0_rd_data_2262;	// matmul/matmul-hw.mlir:20628:36, :20774:5
  //PROBE: c_prev_i_k_4_i_j_11	// matmul/matmul-hw.mlir:20775:5
  assign tk_i_k_4_i_j_11 = _T_2874;	// matmul/matmul-hw.mlir:20777:5
  //PROBE: tk_i_k_4_i_j_11	// matmul/matmul-hw.mlir:20778:5
  wire [31:0] _T_3722 = mult_inst180_result + C_reg_bank4_p0_rd_data_2262;	// matmul/matmul-hw.mlir:20628:36, :20765:28, :20779:13
  assign c_i_k_4_i_j_11 = _T_3722;	// matmul/matmul-hw.mlir:20781:5
  //PROBE: c_i_k_4_i_j_11	// matmul/matmul-hw.mlir:20782:5
  assign _T_408 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20783:13
  assign _T_407 = _T_2902 ? _T_3722 : 32'bx;	// matmul/matmul-hw.mlir:8442:18, :20784:13
  localparam [3:0] _T_3724 = 4'h0;	// matmul/matmul-hw.mlir:20787:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20788:5
    if (rst)	// matmul/matmul-hw.mlir:20788:5
      i_k_next_3723 <= _T_3724;	// matmul/matmul-hw.mlir:20791:7
    else	// matmul/matmul-hw.mlir:20788:5
      i_k_next_3723 <= i_k_next_3720;	// matmul/matmul-hw.mlir:20756:13, :20789:7
  end // always @(posedge)
  assign _T_406 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20793:13
  assign _T_405 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20794:13
  mult mult_inst181 (	// matmul/matmul-hw.mlir:20795:28
    .a      (A_reg_bank181_p0_rd_data),	// matmul/matmul-hw.mlir:12396:33
    .b      (_T_2545),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst181_result)
  );
  assign _T_404 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20796:13
  assign a_i_k_5_i_j_11 = A_reg_bank181_p0_rd_data;	// matmul/matmul-hw.mlir:12396:33, :20798:5
  //PROBE: a_i_k_5_i_j_11	// matmul/matmul-hw.mlir:20799:5
  assign b_i_k_5_i_j_11 = _T_2545;	// matmul/matmul-hw.mlir:20801:5
  //PROBE: b_i_k_5_i_j_11	// matmul/matmul-hw.mlir:20802:5
  assign c_prev_i_k_5_i_j_11 = C_reg_bank5_p0_rd_data_2261;	// matmul/matmul-hw.mlir:20629:36, :20804:5
  //PROBE: c_prev_i_k_5_i_j_11	// matmul/matmul-hw.mlir:20805:5
  assign tk_i_k_5_i_j_11 = _T_2885;	// matmul/matmul-hw.mlir:20807:5
  //PROBE: tk_i_k_5_i_j_11	// matmul/matmul-hw.mlir:20808:5
  wire [31:0] _T_3725 = mult_inst181_result + C_reg_bank5_p0_rd_data_2261;	// matmul/matmul-hw.mlir:20629:36, :20795:28, :20809:13
  assign c_i_k_5_i_j_11 = _T_3725;	// matmul/matmul-hw.mlir:20811:5
  //PROBE: c_i_k_5_i_j_11	// matmul/matmul-hw.mlir:20812:5
  assign _T_403 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20813:13
  assign _T_402 = _T_2907 ? _T_3725 : 32'bx;	// matmul/matmul-hw.mlir:8437:18, :20814:13
  localparam [3:0] _T_3727 = 4'h0;	// matmul/matmul-hw.mlir:20817:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20818:5
    if (rst)	// matmul/matmul-hw.mlir:20818:5
      i_k_next_3726 <= _T_3727;	// matmul/matmul-hw.mlir:20821:7
    else	// matmul/matmul-hw.mlir:20818:5
      i_k_next_3726 <= i_k_next_3723;	// matmul/matmul-hw.mlir:20786:13, :20819:7
  end // always @(posedge)
  assign _T_401 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20823:13
  assign _T_400 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20824:13
  mult mult_inst182 (	// matmul/matmul-hw.mlir:20825:28
    .a      (A_reg_bank182_p0_rd_data),	// matmul/matmul-hw.mlir:12397:33
    .b      (_T_2561),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst182_result)
  );
  assign _T_399 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20826:13
  assign a_i_k_6_i_j_11 = A_reg_bank182_p0_rd_data;	// matmul/matmul-hw.mlir:12397:33, :20828:5
  //PROBE: a_i_k_6_i_j_11	// matmul/matmul-hw.mlir:20829:5
  assign b_i_k_6_i_j_11 = _T_2561;	// matmul/matmul-hw.mlir:20831:5
  //PROBE: b_i_k_6_i_j_11	// matmul/matmul-hw.mlir:20832:5
  assign c_prev_i_k_6_i_j_11 = C_reg_bank6_p0_rd_data_2260;	// matmul/matmul-hw.mlir:20630:36, :20834:5
  //PROBE: c_prev_i_k_6_i_j_11	// matmul/matmul-hw.mlir:20835:5
  assign tk_i_k_6_i_j_11 = _T_2892;	// matmul/matmul-hw.mlir:20837:5
  //PROBE: tk_i_k_6_i_j_11	// matmul/matmul-hw.mlir:20838:5
  wire [31:0] _T_3728 = mult_inst182_result + C_reg_bank6_p0_rd_data_2260;	// matmul/matmul-hw.mlir:20630:36, :20825:28, :20839:13
  assign c_i_k_6_i_j_11 = _T_3728;	// matmul/matmul-hw.mlir:20841:5
  //PROBE: c_i_k_6_i_j_11	// matmul/matmul-hw.mlir:20842:5
  assign _T_398 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20843:13
  assign _T_397 = _T_2912 ? _T_3728 : 32'bx;	// matmul/matmul-hw.mlir:8432:18, :20844:13
  localparam [3:0] _T_3730 = 4'h0;	// matmul/matmul-hw.mlir:20847:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20848:5
    if (rst)	// matmul/matmul-hw.mlir:20848:5
      i_k_next_3729 <= _T_3730;	// matmul/matmul-hw.mlir:20851:7
    else	// matmul/matmul-hw.mlir:20848:5
      i_k_next_3729 <= i_k_next_3726;	// matmul/matmul-hw.mlir:20816:13, :20849:7
  end // always @(posedge)
  assign _T_396 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20853:13
  assign _T_395 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20854:13
  mult mult_inst183 (	// matmul/matmul-hw.mlir:20855:28
    .a      (A_reg_bank183_p0_rd_data),	// matmul/matmul-hw.mlir:12398:33
    .b      (_T_2577),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst183_result)
  );
  assign _T_394 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20856:13
  assign a_i_k_7_i_j_11 = A_reg_bank183_p0_rd_data;	// matmul/matmul-hw.mlir:12398:33, :20858:5
  //PROBE: a_i_k_7_i_j_11	// matmul/matmul-hw.mlir:20859:5
  assign b_i_k_7_i_j_11 = _T_2577;	// matmul/matmul-hw.mlir:20861:5
  //PROBE: b_i_k_7_i_j_11	// matmul/matmul-hw.mlir:20862:5
  assign c_prev_i_k_7_i_j_11 = C_reg_bank7_p0_rd_data_2259;	// matmul/matmul-hw.mlir:20631:36, :20864:5
  //PROBE: c_prev_i_k_7_i_j_11	// matmul/matmul-hw.mlir:20865:5
  assign tk_i_k_7_i_j_11 = _T_2897;	// matmul/matmul-hw.mlir:20867:5
  //PROBE: tk_i_k_7_i_j_11	// matmul/matmul-hw.mlir:20868:5
  wire [31:0] _T_3731 = mult_inst183_result + C_reg_bank7_p0_rd_data_2259;	// matmul/matmul-hw.mlir:20631:36, :20855:28, :20869:13
  assign c_i_k_7_i_j_11 = _T_3731;	// matmul/matmul-hw.mlir:20871:5
  //PROBE: c_i_k_7_i_j_11	// matmul/matmul-hw.mlir:20872:5
  assign _T_393 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20873:13
  assign _T_392 = _T_2917 ? _T_3731 : 32'bx;	// matmul/matmul-hw.mlir:8427:18, :20874:13
  localparam [3:0] _T_3733 = 4'h0;	// matmul/matmul-hw.mlir:20877:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20878:5
    if (rst)	// matmul/matmul-hw.mlir:20878:5
      i_k_next_3732 <= _T_3733;	// matmul/matmul-hw.mlir:20881:7
    else	// matmul/matmul-hw.mlir:20878:5
      i_k_next_3732 <= i_k_next_3729;	// matmul/matmul-hw.mlir:20846:13, :20879:7
  end // always @(posedge)
  assign _T_391 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20883:13
  assign _T_390 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20884:13
  mult mult_inst184 (	// matmul/matmul-hw.mlir:20885:28
    .a      (A_reg_bank184_p0_rd_data),	// matmul/matmul-hw.mlir:12399:33
    .b      (_T_2593),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst184_result)
  );
  assign _T_389 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20886:13
  assign a_i_k_8_i_j_11 = A_reg_bank184_p0_rd_data;	// matmul/matmul-hw.mlir:12399:33, :20888:5
  //PROBE: a_i_k_8_i_j_11	// matmul/matmul-hw.mlir:20889:5
  assign b_i_k_8_i_j_11 = _T_2593;	// matmul/matmul-hw.mlir:20891:5
  //PROBE: b_i_k_8_i_j_11	// matmul/matmul-hw.mlir:20892:5
  assign c_prev_i_k_8_i_j_11 = C_reg_bank8_p0_rd_data_2258;	// matmul/matmul-hw.mlir:20632:36, :20894:5
  //PROBE: c_prev_i_k_8_i_j_11	// matmul/matmul-hw.mlir:20895:5
  assign tk_i_k_8_i_j_11 = _T_2902;	// matmul/matmul-hw.mlir:20897:5
  //PROBE: tk_i_k_8_i_j_11	// matmul/matmul-hw.mlir:20898:5
  wire [31:0] _T_3734 = mult_inst184_result + C_reg_bank8_p0_rd_data_2258;	// matmul/matmul-hw.mlir:20632:36, :20885:28, :20899:13
  assign c_i_k_8_i_j_11 = _T_3734;	// matmul/matmul-hw.mlir:20901:5
  //PROBE: c_i_k_8_i_j_11	// matmul/matmul-hw.mlir:20902:5
  assign _T_388 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20903:13
  assign _T_387 = _T_2922 ? _T_3734 : 32'bx;	// matmul/matmul-hw.mlir:8422:18, :20904:13
  localparam [3:0] _T_3736 = 4'h0;	// matmul/matmul-hw.mlir:20907:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20908:5
    if (rst)	// matmul/matmul-hw.mlir:20908:5
      i_k_next_3735 <= _T_3736;	// matmul/matmul-hw.mlir:20911:7
    else	// matmul/matmul-hw.mlir:20908:5
      i_k_next_3735 <= i_k_next_3732;	// matmul/matmul-hw.mlir:20876:13, :20909:7
  end // always @(posedge)
  assign _T_386 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20913:13
  assign _T_385 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20914:13
  mult mult_inst185 (	// matmul/matmul-hw.mlir:20915:28
    .a      (A_reg_bank185_p0_rd_data),	// matmul/matmul-hw.mlir:12400:33
    .b      (_T_2609),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst185_result)
  );
  assign _T_384 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20916:13
  assign a_i_k_9_i_j_11 = A_reg_bank185_p0_rd_data;	// matmul/matmul-hw.mlir:12400:33, :20918:5
  //PROBE: a_i_k_9_i_j_11	// matmul/matmul-hw.mlir:20919:5
  assign b_i_k_9_i_j_11 = _T_2609;	// matmul/matmul-hw.mlir:20921:5
  //PROBE: b_i_k_9_i_j_11	// matmul/matmul-hw.mlir:20922:5
  assign c_prev_i_k_9_i_j_11 = C_reg_bank9_p0_rd_data_2257;	// matmul/matmul-hw.mlir:20633:36, :20924:5
  //PROBE: c_prev_i_k_9_i_j_11	// matmul/matmul-hw.mlir:20925:5
  assign tk_i_k_9_i_j_11 = _T_2907;	// matmul/matmul-hw.mlir:20927:5
  //PROBE: tk_i_k_9_i_j_11	// matmul/matmul-hw.mlir:20928:5
  wire [31:0] _T_3737 = mult_inst185_result + C_reg_bank9_p0_rd_data_2257;	// matmul/matmul-hw.mlir:20633:36, :20915:28, :20929:13
  assign c_i_k_9_i_j_11 = _T_3737;	// matmul/matmul-hw.mlir:20931:5
  //PROBE: c_i_k_9_i_j_11	// matmul/matmul-hw.mlir:20932:5
  assign _T_383 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20933:13
  assign _T_382 = _T_2927 ? _T_3737 : 32'bx;	// matmul/matmul-hw.mlir:8417:18, :20934:13
  localparam [3:0] _T_3739 = 4'h0;	// matmul/matmul-hw.mlir:20937:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20938:5
    if (rst)	// matmul/matmul-hw.mlir:20938:5
      i_k_next_3738 <= _T_3739;	// matmul/matmul-hw.mlir:20941:7
    else	// matmul/matmul-hw.mlir:20938:5
      i_k_next_3738 <= i_k_next_3735;	// matmul/matmul-hw.mlir:20906:13, :20939:7
  end // always @(posedge)
  assign _T_381 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20943:13
  assign _T_380 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20944:13
  mult mult_inst186 (	// matmul/matmul-hw.mlir:20945:28
    .a      (A_reg_bank186_p0_rd_data),	// matmul/matmul-hw.mlir:12401:33
    .b      (_T_2625),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst186_result)
  );
  assign _T_379 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20946:13
  assign a_i_k_10_i_j_11 = A_reg_bank186_p0_rd_data;	// matmul/matmul-hw.mlir:12401:33, :20948:5
  //PROBE: a_i_k_10_i_j_11	// matmul/matmul-hw.mlir:20949:5
  assign b_i_k_10_i_j_11 = _T_2625;	// matmul/matmul-hw.mlir:20951:5
  //PROBE: b_i_k_10_i_j_11	// matmul/matmul-hw.mlir:20952:5
  assign c_prev_i_k_10_i_j_11 = C_reg_bank10_p0_rd_data_2256;	// matmul/matmul-hw.mlir:20634:37, :20954:5
  //PROBE: c_prev_i_k_10_i_j_11	// matmul/matmul-hw.mlir:20955:5
  assign tk_i_k_10_i_j_11 = _T_2912;	// matmul/matmul-hw.mlir:20957:5
  //PROBE: tk_i_k_10_i_j_11	// matmul/matmul-hw.mlir:20958:5
  wire [31:0] _T_3740 = mult_inst186_result + C_reg_bank10_p0_rd_data_2256;	// matmul/matmul-hw.mlir:20634:37, :20945:28, :20959:13
  assign c_i_k_10_i_j_11 = _T_3740;	// matmul/matmul-hw.mlir:20961:5
  //PROBE: c_i_k_10_i_j_11	// matmul/matmul-hw.mlir:20962:5
  assign _T_378 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20963:13
  assign _T_377 = _T_2932 ? _T_3740 : 32'bx;	// matmul/matmul-hw.mlir:8412:18, :20964:13
  localparam [3:0] _T_3742 = 4'h0;	// matmul/matmul-hw.mlir:20967:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20968:5
    if (rst)	// matmul/matmul-hw.mlir:20968:5
      i_k_next_3741 <= _T_3742;	// matmul/matmul-hw.mlir:20971:7
    else	// matmul/matmul-hw.mlir:20968:5
      i_k_next_3741 <= i_k_next_3738;	// matmul/matmul-hw.mlir:20936:13, :20969:7
  end // always @(posedge)
  assign _T_376 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20973:13
  assign _T_375 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20974:13
  mult mult_inst187 (	// matmul/matmul-hw.mlir:20975:28
    .a      (A_reg_bank187_p0_rd_data),	// matmul/matmul-hw.mlir:12402:33
    .b      (_T_2641),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst187_result)
  );
  assign _T_374 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20976:13
  assign a_i_k_11_i_j_11 = A_reg_bank187_p0_rd_data;	// matmul/matmul-hw.mlir:12402:33, :20978:5
  //PROBE: a_i_k_11_i_j_11	// matmul/matmul-hw.mlir:20979:5
  assign b_i_k_11_i_j_11 = _T_2641;	// matmul/matmul-hw.mlir:20981:5
  //PROBE: b_i_k_11_i_j_11	// matmul/matmul-hw.mlir:20982:5
  assign c_prev_i_k_11_i_j_11 = C_reg_bank11_p0_rd_data_2255;	// matmul/matmul-hw.mlir:20635:37, :20984:5
  //PROBE: c_prev_i_k_11_i_j_11	// matmul/matmul-hw.mlir:20985:5
  assign tk_i_k_11_i_j_11 = _T_2917;	// matmul/matmul-hw.mlir:20987:5
  //PROBE: tk_i_k_11_i_j_11	// matmul/matmul-hw.mlir:20988:5
  wire [31:0] _T_3743 = mult_inst187_result + C_reg_bank11_p0_rd_data_2255;	// matmul/matmul-hw.mlir:20635:37, :20975:28, :20989:13
  assign c_i_k_11_i_j_11 = _T_3743;	// matmul/matmul-hw.mlir:20991:5
  //PROBE: c_i_k_11_i_j_11	// matmul/matmul-hw.mlir:20992:5
  assign _T_373 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :20993:13
  assign _T_372 = _T_2937 ? _T_3743 : 32'bx;	// matmul/matmul-hw.mlir:8407:18, :20994:13
  localparam [3:0] _T_3745 = 4'h0;	// matmul/matmul-hw.mlir:20997:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:20998:5
    if (rst)	// matmul/matmul-hw.mlir:20998:5
      i_k_next_3744 <= _T_3745;	// matmul/matmul-hw.mlir:21001:7
    else	// matmul/matmul-hw.mlir:20998:5
      i_k_next_3744 <= i_k_next_3741;	// matmul/matmul-hw.mlir:20966:13, :20999:7
  end // always @(posedge)
  assign _T_371 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21003:13
  assign _T_370 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21004:13
  mult mult_inst188 (	// matmul/matmul-hw.mlir:21005:28
    .a      (A_reg_bank188_p0_rd_data),	// matmul/matmul-hw.mlir:12403:33
    .b      (_T_2657),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst188_result)
  );
  assign _T_369 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21006:13
  assign a_i_k_12_i_j_11 = A_reg_bank188_p0_rd_data;	// matmul/matmul-hw.mlir:12403:33, :21008:5
  //PROBE: a_i_k_12_i_j_11	// matmul/matmul-hw.mlir:21009:5
  assign b_i_k_12_i_j_11 = _T_2657;	// matmul/matmul-hw.mlir:21011:5
  //PROBE: b_i_k_12_i_j_11	// matmul/matmul-hw.mlir:21012:5
  assign c_prev_i_k_12_i_j_11 = C_reg_bank12_p0_rd_data_2254;	// matmul/matmul-hw.mlir:20636:37, :21014:5
  //PROBE: c_prev_i_k_12_i_j_11	// matmul/matmul-hw.mlir:21015:5
  assign tk_i_k_12_i_j_11 = _T_2922;	// matmul/matmul-hw.mlir:21017:5
  //PROBE: tk_i_k_12_i_j_11	// matmul/matmul-hw.mlir:21018:5
  wire [31:0] _T_3746 = mult_inst188_result + C_reg_bank12_p0_rd_data_2254;	// matmul/matmul-hw.mlir:20636:37, :21005:28, :21019:13
  assign c_i_k_12_i_j_11 = _T_3746;	// matmul/matmul-hw.mlir:21021:5
  //PROBE: c_i_k_12_i_j_11	// matmul/matmul-hw.mlir:21022:5
  assign _T_368 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21023:13
  assign _T_367 = _T_2942 ? _T_3746 : 32'bx;	// matmul/matmul-hw.mlir:8402:18, :21024:13
  localparam [3:0] _T_3748 = 4'h0;	// matmul/matmul-hw.mlir:21027:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21028:5
    if (rst)	// matmul/matmul-hw.mlir:21028:5
      i_k_next_3747 <= _T_3748;	// matmul/matmul-hw.mlir:21031:7
    else	// matmul/matmul-hw.mlir:21028:5
      i_k_next_3747 <= i_k_next_3744;	// matmul/matmul-hw.mlir:20996:13, :21029:7
  end // always @(posedge)
  assign _T_366 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21033:13
  assign _T_365 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21034:13
  mult mult_inst189 (	// matmul/matmul-hw.mlir:21035:28
    .a      (A_reg_bank189_p0_rd_data),	// matmul/matmul-hw.mlir:12404:33
    .b      (_T_2673),
    .t      (_T_2937),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst189_result)
  );
  assign _T_364 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21036:13
  assign a_i_k_13_i_j_11 = A_reg_bank189_p0_rd_data;	// matmul/matmul-hw.mlir:12404:33, :21038:5
  //PROBE: a_i_k_13_i_j_11	// matmul/matmul-hw.mlir:21039:5
  assign b_i_k_13_i_j_11 = _T_2673;	// matmul/matmul-hw.mlir:21041:5
  //PROBE: b_i_k_13_i_j_11	// matmul/matmul-hw.mlir:21042:5
  assign c_prev_i_k_13_i_j_11 = C_reg_bank13_p0_rd_data_2253;	// matmul/matmul-hw.mlir:20637:37, :21044:5
  //PROBE: c_prev_i_k_13_i_j_11	// matmul/matmul-hw.mlir:21045:5
  assign tk_i_k_13_i_j_11 = _T_2927;	// matmul/matmul-hw.mlir:21047:5
  //PROBE: tk_i_k_13_i_j_11	// matmul/matmul-hw.mlir:21048:5
  wire [31:0] _T_3749 = mult_inst189_result + C_reg_bank13_p0_rd_data_2253;	// matmul/matmul-hw.mlir:20637:37, :21035:28, :21049:13
  assign c_i_k_13_i_j_11 = _T_3749;	// matmul/matmul-hw.mlir:21051:5
  //PROBE: c_i_k_13_i_j_11	// matmul/matmul-hw.mlir:21052:5
  assign _T_363 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21053:13
  assign _T_362 = _T_2947 ? _T_3749 : 32'bx;	// matmul/matmul-hw.mlir:8397:18, :21054:13
  localparam [3:0] _T_3751 = 4'h0;	// matmul/matmul-hw.mlir:21057:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21058:5
    if (rst)	// matmul/matmul-hw.mlir:21058:5
      i_k_next_3750 <= _T_3751;	// matmul/matmul-hw.mlir:21061:7
    else	// matmul/matmul-hw.mlir:21058:5
      i_k_next_3750 <= i_k_next_3747;	// matmul/matmul-hw.mlir:21026:13, :21059:7
  end // always @(posedge)
  assign _T_361 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21063:13
  assign _T_360 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21064:13
  mult mult_inst190 (	// matmul/matmul-hw.mlir:21065:28
    .a      (A_reg_bank190_p0_rd_data),	// matmul/matmul-hw.mlir:12405:33
    .b      (_T_2689),
    .t      (_T_2942),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst190_result)
  );
  assign _T_359 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21066:13
  assign a_i_k_14_i_j_11 = A_reg_bank190_p0_rd_data;	// matmul/matmul-hw.mlir:12405:33, :21068:5
  //PROBE: a_i_k_14_i_j_11	// matmul/matmul-hw.mlir:21069:5
  assign b_i_k_14_i_j_11 = _T_2689;	// matmul/matmul-hw.mlir:21071:5
  //PROBE: b_i_k_14_i_j_11	// matmul/matmul-hw.mlir:21072:5
  assign c_prev_i_k_14_i_j_11 = C_reg_bank14_p0_rd_data_2252;	// matmul/matmul-hw.mlir:20638:37, :21074:5
  //PROBE: c_prev_i_k_14_i_j_11	// matmul/matmul-hw.mlir:21075:5
  assign tk_i_k_14_i_j_11 = _T_2932;	// matmul/matmul-hw.mlir:21077:5
  //PROBE: tk_i_k_14_i_j_11	// matmul/matmul-hw.mlir:21078:5
  wire [31:0] _T_3752 = mult_inst190_result + C_reg_bank14_p0_rd_data_2252;	// matmul/matmul-hw.mlir:20638:37, :21065:28, :21079:13
  assign c_i_k_14_i_j_11 = _T_3752;	// matmul/matmul-hw.mlir:21081:5
  //PROBE: c_i_k_14_i_j_11	// matmul/matmul-hw.mlir:21082:5
  assign _T_358 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21083:13
  assign _T_357 = _T_2952 ? _T_3752 : 32'bx;	// matmul/matmul-hw.mlir:8392:18, :21084:13
  localparam [3:0] _T_3754 = 4'h0;	// matmul/matmul-hw.mlir:21087:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21088:5
    if (rst)	// matmul/matmul-hw.mlir:21088:5
      i_k_next_3753 <= _T_3754;	// matmul/matmul-hw.mlir:21091:7
    else	// matmul/matmul-hw.mlir:21088:5
      i_k_next_3753 <= i_k_next_3750;	// matmul/matmul-hw.mlir:21056:13, :21089:7
  end // always @(posedge)
  assign _T_356 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21093:13
  assign _T_355 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21094:13
  mult mult_inst191 (	// matmul/matmul-hw.mlir:21095:28
    .a      (A_reg_bank191_p0_rd_data),	// matmul/matmul-hw.mlir:12406:33
    .b      (_T_2705),
    .t      (_T_2947),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst191_result)
  );
  assign _T_354 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21096:13
  assign a_i_k_15_i_j_11 = A_reg_bank191_p0_rd_data;	// matmul/matmul-hw.mlir:12406:33, :21098:5
  //PROBE: a_i_k_15_i_j_11	// matmul/matmul-hw.mlir:21099:5
  assign b_i_k_15_i_j_11 = _T_2705;	// matmul/matmul-hw.mlir:21101:5
  //PROBE: b_i_k_15_i_j_11	// matmul/matmul-hw.mlir:21102:5
  assign c_prev_i_k_15_i_j_11 = C_reg_bank15_p0_rd_data_2251;	// matmul/matmul-hw.mlir:20639:37, :21104:5
  //PROBE: c_prev_i_k_15_i_j_11	// matmul/matmul-hw.mlir:21105:5
  assign tk_i_k_15_i_j_11 = _T_2937;	// matmul/matmul-hw.mlir:21107:5
  //PROBE: tk_i_k_15_i_j_11	// matmul/matmul-hw.mlir:21108:5
  wire [31:0] _T_3755 = mult_inst191_result + C_reg_bank15_p0_rd_data_2251;	// matmul/matmul-hw.mlir:20639:37, :21095:28, :21109:13
  assign c_i_k_15_i_j_11 = _T_3755;	// matmul/matmul-hw.mlir:21111:5
  //PROBE: c_i_k_15_i_j_11	// matmul/matmul-hw.mlir:21112:5
  assign _T_353 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21113:13
  assign _T_352 = _T_2957 ? _T_3755 : 32'bx;	// matmul/matmul-hw.mlir:8387:18, :21114:13
  localparam [3:0] _T_3757 = 4'h0;	// matmul/matmul-hw.mlir:21117:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21118:5
    if (rst)	// matmul/matmul-hw.mlir:21118:5
      i_k_next_3756 <= _T_3757;	// matmul/matmul-hw.mlir:21121:7
    else	// matmul/matmul-hw.mlir:21118:5
      i_k_next_3756 <= i_k_next_3753;	// matmul/matmul-hw.mlir:21086:13, :21119:7
  end // always @(posedge)
  assign _T_351 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21123:13
  wire [3:0][3:0] _T_3759 = i_delayed_3758;	// matmul/matmul-hw.mlir:21125:13
  wire [3:0][3:0] _T_3760 = {_T_3759[2'h0+:3], {{i_k_next_3756}}};	// matmul/matmul-hw.mlir:21116:13, :21126:19, :21127:13, :21128:13, :21129:13
  wire [3:0][3:0] _T_3761 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:21130:19, :21131:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21132:5
    if (rst)	// matmul/matmul-hw.mlir:21132:5
      i_delayed_3758 <= _T_3761;	// matmul/matmul-hw.mlir:21135:7
    else	// matmul/matmul-hw.mlir:21132:5
      i_delayed_3758 <= _T_3760;	// matmul/matmul-hw.mlir:21133:7
  end // always @(posedge)
  assign _T_350 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21139:13
  assign _T_349 = _T_2962 ? i_delayed_3758[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8384:17, :21125:13, :21137:20, :21138:13, :21140:13
  assign _T_348 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21141:13
  assign _T_347 = _T_2962 ? C_reg_bank16_p0_rd_data_2250 : 32'bx;	// matmul/matmul-hw.mlir:8382:18, :20640:37, :21142:13
  localparam [3:0] _T_3763 = 4'h0;	// matmul/matmul-hw.mlir:21145:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21146:5
    if (rst)	// matmul/matmul-hw.mlir:21146:5
      i_j_next_3762 <= _T_3763;	// matmul/matmul-hw.mlir:21149:7
    else	// matmul/matmul-hw.mlir:21146:5
      i_j_next_3762 <= i_j_next_3691;	// matmul/matmul-hw.mlir:20549:13, :21147:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3764 (	// matmul/matmul-hw.mlir:21219:36
    .p0_rd_en   (_T_342),	// matmul/matmul-hw.mlir:21241:13
    .p1_wr_en   (_T_346),	// matmul/matmul-hw.mlir:21236:13
    .p1_wr_data (_T_345),	// matmul/matmul-hw.mlir:21237:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2249)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3765 (	// matmul/matmul-hw.mlir:21220:36
    .p0_rd_en   (_T_337),	// matmul/matmul-hw.mlir:21271:13
    .p1_wr_en   (_T_341),	// matmul/matmul-hw.mlir:21258:13
    .p1_wr_data (_T_340),	// matmul/matmul-hw.mlir:21259:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2248)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3766 (	// matmul/matmul-hw.mlir:21221:36
    .p0_rd_en   (_T_332),	// matmul/matmul-hw.mlir:21301:13
    .p1_wr_en   (_T_336),	// matmul/matmul-hw.mlir:21288:13
    .p1_wr_data (_T_335),	// matmul/matmul-hw.mlir:21289:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2247)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3767 (	// matmul/matmul-hw.mlir:21222:36
    .p0_rd_en   (_T_327),	// matmul/matmul-hw.mlir:21331:13
    .p1_wr_en   (_T_331),	// matmul/matmul-hw.mlir:21318:13
    .p1_wr_data (_T_330),	// matmul/matmul-hw.mlir:21319:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2246)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3768 (	// matmul/matmul-hw.mlir:21223:36
    .p0_rd_en   (_T_322),	// matmul/matmul-hw.mlir:21361:13
    .p1_wr_en   (_T_326),	// matmul/matmul-hw.mlir:21348:13
    .p1_wr_data (_T_325),	// matmul/matmul-hw.mlir:21349:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2245)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3769 (	// matmul/matmul-hw.mlir:21224:36
    .p0_rd_en   (_T_317),	// matmul/matmul-hw.mlir:21391:13
    .p1_wr_en   (_T_321),	// matmul/matmul-hw.mlir:21378:13
    .p1_wr_data (_T_320),	// matmul/matmul-hw.mlir:21379:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2244)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3770 (	// matmul/matmul-hw.mlir:21225:36
    .p0_rd_en   (_T_312),	// matmul/matmul-hw.mlir:21421:13
    .p1_wr_en   (_T_316),	// matmul/matmul-hw.mlir:21408:13
    .p1_wr_data (_T_315),	// matmul/matmul-hw.mlir:21409:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2243)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3771 (	// matmul/matmul-hw.mlir:21226:36
    .p0_rd_en   (_T_307),	// matmul/matmul-hw.mlir:21451:13
    .p1_wr_en   (_T_311),	// matmul/matmul-hw.mlir:21438:13
    .p1_wr_data (_T_310),	// matmul/matmul-hw.mlir:21439:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2242)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3772 (	// matmul/matmul-hw.mlir:21227:36
    .p0_rd_en   (_T_302),	// matmul/matmul-hw.mlir:21481:13
    .p1_wr_en   (_T_306),	// matmul/matmul-hw.mlir:21468:13
    .p1_wr_data (_T_305),	// matmul/matmul-hw.mlir:21469:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2241)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3773 (	// matmul/matmul-hw.mlir:21228:36
    .p0_rd_en   (_T_297),	// matmul/matmul-hw.mlir:21511:13
    .p1_wr_en   (_T_301),	// matmul/matmul-hw.mlir:21498:13
    .p1_wr_data (_T_300),	// matmul/matmul-hw.mlir:21499:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2240)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3774 (	// matmul/matmul-hw.mlir:21229:37
    .p0_rd_en   (_T_292),	// matmul/matmul-hw.mlir:21541:13
    .p1_wr_en   (_T_296),	// matmul/matmul-hw.mlir:21528:13
    .p1_wr_data (_T_295),	// matmul/matmul-hw.mlir:21529:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2239)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3775 (	// matmul/matmul-hw.mlir:21230:37
    .p0_rd_en   (_T_287),	// matmul/matmul-hw.mlir:21571:13
    .p1_wr_en   (_T_291),	// matmul/matmul-hw.mlir:21558:13
    .p1_wr_data (_T_290),	// matmul/matmul-hw.mlir:21559:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2238)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3776 (	// matmul/matmul-hw.mlir:21231:37
    .p0_rd_en   (_T_282),	// matmul/matmul-hw.mlir:21601:13
    .p1_wr_en   (_T_286),	// matmul/matmul-hw.mlir:21588:13
    .p1_wr_data (_T_285),	// matmul/matmul-hw.mlir:21589:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2237)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3777 (	// matmul/matmul-hw.mlir:21232:37
    .p0_rd_en   (_T_277),	// matmul/matmul-hw.mlir:21631:13
    .p1_wr_en   (_T_281),	// matmul/matmul-hw.mlir:21618:13
    .p1_wr_data (_T_280),	// matmul/matmul-hw.mlir:21619:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2236)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3778 (	// matmul/matmul-hw.mlir:21233:37
    .p0_rd_en   (_T_272),	// matmul/matmul-hw.mlir:21661:13
    .p1_wr_en   (_T_276),	// matmul/matmul-hw.mlir:21648:13
    .p1_wr_data (_T_275),	// matmul/matmul-hw.mlir:21649:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2235)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3779 (	// matmul/matmul-hw.mlir:21234:37
    .p0_rd_en   (_T_267),	// matmul/matmul-hw.mlir:21691:13
    .p1_wr_en   (_T_271),	// matmul/matmul-hw.mlir:21678:13
    .p1_wr_data (_T_270),	// matmul/matmul-hw.mlir:21679:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2234)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3780 (	// matmul/matmul-hw.mlir:21235:37
    .p0_rd_en   (_T_264),	// matmul/matmul-hw.mlir:21733:13
    .p1_wr_en   (_T_266),	// matmul/matmul-hw.mlir:21708:13
    .p1_wr_data (_T_265),	// matmul/matmul-hw.mlir:21709:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2233)
  );
  assign _T_346 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21236:13
  assign _T_345 = _T_2874 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8380:18, :21237:13
  assign _T_344 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21238:13
  assign _T_343 = _T_2863 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21239:13
  mult mult_inst192 (	// matmul/matmul-hw.mlir:21240:28
    .a      (A_reg_bank192_p0_rd_data),	// matmul/matmul-hw.mlir:12407:33
    .b      (_T_2466),
    .t      (_T_2863),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst192_result)
  );
  assign _T_342 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21241:13
  assign a_i_k_0_i_j_12 = A_reg_bank192_p0_rd_data;	// matmul/matmul-hw.mlir:12407:33, :21243:5
  //PROBE: a_i_k_0_i_j_12	// matmul/matmul-hw.mlir:21244:5
  assign b_i_k_0_i_j_12 = _T_2466;	// matmul/matmul-hw.mlir:21246:5
  //PROBE: b_i_k_0_i_j_12	// matmul/matmul-hw.mlir:21247:5
  assign c_prev_i_k_0_i_j_12 = C_reg_bank0_p0_rd_data_2249;	// matmul/matmul-hw.mlir:21219:36, :21249:5
  //PROBE: c_prev_i_k_0_i_j_12	// matmul/matmul-hw.mlir:21250:5
  assign tk_i_k_0_i_j_12 = _T_2841;	// matmul/matmul-hw.mlir:21252:5
  //PROBE: tk_i_k_0_i_j_12	// matmul/matmul-hw.mlir:21253:5
  wire [31:0] _T_3781 = mult_inst192_result + C_reg_bank0_p0_rd_data_2249;	// matmul/matmul-hw.mlir:21219:36, :21240:28, :21254:13
  assign c_i_k_0_i_j_12 = _T_3781;	// matmul/matmul-hw.mlir:21256:5
  //PROBE: c_i_k_0_i_j_12	// matmul/matmul-hw.mlir:21257:5
  assign _T_341 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21258:13
  assign _T_340 = _T_2885 ? _T_3781 : 32'bx;	// matmul/matmul-hw.mlir:8375:18, :21259:13
  localparam [3:0] _T_3783 = 4'h0;	// matmul/matmul-hw.mlir:21262:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21263:5
    if (rst)	// matmul/matmul-hw.mlir:21263:5
      i_k_next_3782 <= _T_3783;	// matmul/matmul-hw.mlir:21266:7
    else	// matmul/matmul-hw.mlir:21263:5
      i_k_next_3782 <= i_j_next_3762;	// matmul/matmul-hw.mlir:21144:13, :21264:7
  end // always @(posedge)
  assign _T_339 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21268:13
  assign _T_338 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21269:13
  mult mult_inst193 (	// matmul/matmul-hw.mlir:21270:28
    .a      (A_reg_bank193_p0_rd_data),	// matmul/matmul-hw.mlir:12408:33
    .b      (_T_2482),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst193_result)
  );
  assign _T_337 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21271:13
  assign a_i_k_1_i_j_12 = A_reg_bank193_p0_rd_data;	// matmul/matmul-hw.mlir:12408:33, :21273:5
  //PROBE: a_i_k_1_i_j_12	// matmul/matmul-hw.mlir:21274:5
  assign b_i_k_1_i_j_12 = _T_2482;	// matmul/matmul-hw.mlir:21276:5
  //PROBE: b_i_k_1_i_j_12	// matmul/matmul-hw.mlir:21277:5
  assign c_prev_i_k_1_i_j_12 = C_reg_bank1_p0_rd_data_2248;	// matmul/matmul-hw.mlir:21220:36, :21279:5
  //PROBE: c_prev_i_k_1_i_j_12	// matmul/matmul-hw.mlir:21280:5
  assign tk_i_k_1_i_j_12 = _T_2852;	// matmul/matmul-hw.mlir:21282:5
  //PROBE: tk_i_k_1_i_j_12	// matmul/matmul-hw.mlir:21283:5
  wire [31:0] _T_3784 = mult_inst193_result + C_reg_bank1_p0_rd_data_2248;	// matmul/matmul-hw.mlir:21220:36, :21270:28, :21284:13
  assign c_i_k_1_i_j_12 = _T_3784;	// matmul/matmul-hw.mlir:21286:5
  //PROBE: c_i_k_1_i_j_12	// matmul/matmul-hw.mlir:21287:5
  assign _T_336 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21288:13
  assign _T_335 = _T_2892 ? _T_3784 : 32'bx;	// matmul/matmul-hw.mlir:8370:18, :21289:13
  localparam [3:0] _T_3786 = 4'h0;	// matmul/matmul-hw.mlir:21292:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21293:5
    if (rst)	// matmul/matmul-hw.mlir:21293:5
      i_k_next_3785 <= _T_3786;	// matmul/matmul-hw.mlir:21296:7
    else	// matmul/matmul-hw.mlir:21293:5
      i_k_next_3785 <= i_k_next_3782;	// matmul/matmul-hw.mlir:21261:13, :21294:7
  end // always @(posedge)
  assign _T_334 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21298:13
  assign _T_333 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21299:13
  mult mult_inst194 (	// matmul/matmul-hw.mlir:21300:28
    .a      (A_reg_bank194_p0_rd_data),	// matmul/matmul-hw.mlir:12409:33
    .b      (_T_2498),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst194_result)
  );
  assign _T_332 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21301:13
  assign a_i_k_2_i_j_12 = A_reg_bank194_p0_rd_data;	// matmul/matmul-hw.mlir:12409:33, :21303:5
  //PROBE: a_i_k_2_i_j_12	// matmul/matmul-hw.mlir:21304:5
  assign b_i_k_2_i_j_12 = _T_2498;	// matmul/matmul-hw.mlir:21306:5
  //PROBE: b_i_k_2_i_j_12	// matmul/matmul-hw.mlir:21307:5
  assign c_prev_i_k_2_i_j_12 = C_reg_bank2_p0_rd_data_2247;	// matmul/matmul-hw.mlir:21221:36, :21309:5
  //PROBE: c_prev_i_k_2_i_j_12	// matmul/matmul-hw.mlir:21310:5
  assign tk_i_k_2_i_j_12 = _T_2863;	// matmul/matmul-hw.mlir:21312:5
  //PROBE: tk_i_k_2_i_j_12	// matmul/matmul-hw.mlir:21313:5
  wire [31:0] _T_3787 = mult_inst194_result + C_reg_bank2_p0_rd_data_2247;	// matmul/matmul-hw.mlir:21221:36, :21300:28, :21314:13
  assign c_i_k_2_i_j_12 = _T_3787;	// matmul/matmul-hw.mlir:21316:5
  //PROBE: c_i_k_2_i_j_12	// matmul/matmul-hw.mlir:21317:5
  assign _T_331 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21318:13
  assign _T_330 = _T_2897 ? _T_3787 : 32'bx;	// matmul/matmul-hw.mlir:8365:18, :21319:13
  localparam [3:0] _T_3789 = 4'h0;	// matmul/matmul-hw.mlir:21322:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21323:5
    if (rst)	// matmul/matmul-hw.mlir:21323:5
      i_k_next_3788 <= _T_3789;	// matmul/matmul-hw.mlir:21326:7
    else	// matmul/matmul-hw.mlir:21323:5
      i_k_next_3788 <= i_k_next_3785;	// matmul/matmul-hw.mlir:21291:13, :21324:7
  end // always @(posedge)
  assign _T_329 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21328:13
  assign _T_328 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21329:13
  mult mult_inst195 (	// matmul/matmul-hw.mlir:21330:28
    .a      (A_reg_bank195_p0_rd_data),	// matmul/matmul-hw.mlir:12410:33
    .b      (_T_2514),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst195_result)
  );
  assign _T_327 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21331:13
  assign a_i_k_3_i_j_12 = A_reg_bank195_p0_rd_data;	// matmul/matmul-hw.mlir:12410:33, :21333:5
  //PROBE: a_i_k_3_i_j_12	// matmul/matmul-hw.mlir:21334:5
  assign b_i_k_3_i_j_12 = _T_2514;	// matmul/matmul-hw.mlir:21336:5
  //PROBE: b_i_k_3_i_j_12	// matmul/matmul-hw.mlir:21337:5
  assign c_prev_i_k_3_i_j_12 = C_reg_bank3_p0_rd_data_2246;	// matmul/matmul-hw.mlir:21222:36, :21339:5
  //PROBE: c_prev_i_k_3_i_j_12	// matmul/matmul-hw.mlir:21340:5
  assign tk_i_k_3_i_j_12 = _T_2874;	// matmul/matmul-hw.mlir:21342:5
  //PROBE: tk_i_k_3_i_j_12	// matmul/matmul-hw.mlir:21343:5
  wire [31:0] _T_3790 = mult_inst195_result + C_reg_bank3_p0_rd_data_2246;	// matmul/matmul-hw.mlir:21222:36, :21330:28, :21344:13
  assign c_i_k_3_i_j_12 = _T_3790;	// matmul/matmul-hw.mlir:21346:5
  //PROBE: c_i_k_3_i_j_12	// matmul/matmul-hw.mlir:21347:5
  assign _T_326 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21348:13
  assign _T_325 = _T_2902 ? _T_3790 : 32'bx;	// matmul/matmul-hw.mlir:8360:18, :21349:13
  localparam [3:0] _T_3792 = 4'h0;	// matmul/matmul-hw.mlir:21352:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21353:5
    if (rst)	// matmul/matmul-hw.mlir:21353:5
      i_k_next_3791 <= _T_3792;	// matmul/matmul-hw.mlir:21356:7
    else	// matmul/matmul-hw.mlir:21353:5
      i_k_next_3791 <= i_k_next_3788;	// matmul/matmul-hw.mlir:21321:13, :21354:7
  end // always @(posedge)
  assign _T_324 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21358:13
  assign _T_323 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21359:13
  mult mult_inst196 (	// matmul/matmul-hw.mlir:21360:28
    .a      (A_reg_bank196_p0_rd_data),	// matmul/matmul-hw.mlir:12411:33
    .b      (_T_2530),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst196_result)
  );
  assign _T_322 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21361:13
  assign a_i_k_4_i_j_12 = A_reg_bank196_p0_rd_data;	// matmul/matmul-hw.mlir:12411:33, :21363:5
  //PROBE: a_i_k_4_i_j_12	// matmul/matmul-hw.mlir:21364:5
  assign b_i_k_4_i_j_12 = _T_2530;	// matmul/matmul-hw.mlir:21366:5
  //PROBE: b_i_k_4_i_j_12	// matmul/matmul-hw.mlir:21367:5
  assign c_prev_i_k_4_i_j_12 = C_reg_bank4_p0_rd_data_2245;	// matmul/matmul-hw.mlir:21223:36, :21369:5
  //PROBE: c_prev_i_k_4_i_j_12	// matmul/matmul-hw.mlir:21370:5
  assign tk_i_k_4_i_j_12 = _T_2885;	// matmul/matmul-hw.mlir:21372:5
  //PROBE: tk_i_k_4_i_j_12	// matmul/matmul-hw.mlir:21373:5
  wire [31:0] _T_3793 = mult_inst196_result + C_reg_bank4_p0_rd_data_2245;	// matmul/matmul-hw.mlir:21223:36, :21360:28, :21374:13
  assign c_i_k_4_i_j_12 = _T_3793;	// matmul/matmul-hw.mlir:21376:5
  //PROBE: c_i_k_4_i_j_12	// matmul/matmul-hw.mlir:21377:5
  assign _T_321 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21378:13
  assign _T_320 = _T_2907 ? _T_3793 : 32'bx;	// matmul/matmul-hw.mlir:8355:18, :21379:13
  localparam [3:0] _T_3795 = 4'h0;	// matmul/matmul-hw.mlir:21382:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21383:5
    if (rst)	// matmul/matmul-hw.mlir:21383:5
      i_k_next_3794 <= _T_3795;	// matmul/matmul-hw.mlir:21386:7
    else	// matmul/matmul-hw.mlir:21383:5
      i_k_next_3794 <= i_k_next_3791;	// matmul/matmul-hw.mlir:21351:13, :21384:7
  end // always @(posedge)
  assign _T_319 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21388:13
  assign _T_318 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21389:13
  mult mult_inst197 (	// matmul/matmul-hw.mlir:21390:28
    .a      (A_reg_bank197_p0_rd_data),	// matmul/matmul-hw.mlir:12412:33
    .b      (_T_2546),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst197_result)
  );
  assign _T_317 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21391:13
  assign a_i_k_5_i_j_12 = A_reg_bank197_p0_rd_data;	// matmul/matmul-hw.mlir:12412:33, :21393:5
  //PROBE: a_i_k_5_i_j_12	// matmul/matmul-hw.mlir:21394:5
  assign b_i_k_5_i_j_12 = _T_2546;	// matmul/matmul-hw.mlir:21396:5
  //PROBE: b_i_k_5_i_j_12	// matmul/matmul-hw.mlir:21397:5
  assign c_prev_i_k_5_i_j_12 = C_reg_bank5_p0_rd_data_2244;	// matmul/matmul-hw.mlir:21224:36, :21399:5
  //PROBE: c_prev_i_k_5_i_j_12	// matmul/matmul-hw.mlir:21400:5
  assign tk_i_k_5_i_j_12 = _T_2892;	// matmul/matmul-hw.mlir:21402:5
  //PROBE: tk_i_k_5_i_j_12	// matmul/matmul-hw.mlir:21403:5
  wire [31:0] _T_3796 = mult_inst197_result + C_reg_bank5_p0_rd_data_2244;	// matmul/matmul-hw.mlir:21224:36, :21390:28, :21404:13
  assign c_i_k_5_i_j_12 = _T_3796;	// matmul/matmul-hw.mlir:21406:5
  //PROBE: c_i_k_5_i_j_12	// matmul/matmul-hw.mlir:21407:5
  assign _T_316 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21408:13
  assign _T_315 = _T_2912 ? _T_3796 : 32'bx;	// matmul/matmul-hw.mlir:8350:18, :21409:13
  localparam [3:0] _T_3798 = 4'h0;	// matmul/matmul-hw.mlir:21412:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21413:5
    if (rst)	// matmul/matmul-hw.mlir:21413:5
      i_k_next_3797 <= _T_3798;	// matmul/matmul-hw.mlir:21416:7
    else	// matmul/matmul-hw.mlir:21413:5
      i_k_next_3797 <= i_k_next_3794;	// matmul/matmul-hw.mlir:21381:13, :21414:7
  end // always @(posedge)
  assign _T_314 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21418:13
  assign _T_313 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21419:13
  mult mult_inst198 (	// matmul/matmul-hw.mlir:21420:28
    .a      (A_reg_bank198_p0_rd_data),	// matmul/matmul-hw.mlir:12413:33
    .b      (_T_2562),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst198_result)
  );
  assign _T_312 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21421:13
  assign a_i_k_6_i_j_12 = A_reg_bank198_p0_rd_data;	// matmul/matmul-hw.mlir:12413:33, :21423:5
  //PROBE: a_i_k_6_i_j_12	// matmul/matmul-hw.mlir:21424:5
  assign b_i_k_6_i_j_12 = _T_2562;	// matmul/matmul-hw.mlir:21426:5
  //PROBE: b_i_k_6_i_j_12	// matmul/matmul-hw.mlir:21427:5
  assign c_prev_i_k_6_i_j_12 = C_reg_bank6_p0_rd_data_2243;	// matmul/matmul-hw.mlir:21225:36, :21429:5
  //PROBE: c_prev_i_k_6_i_j_12	// matmul/matmul-hw.mlir:21430:5
  assign tk_i_k_6_i_j_12 = _T_2897;	// matmul/matmul-hw.mlir:21432:5
  //PROBE: tk_i_k_6_i_j_12	// matmul/matmul-hw.mlir:21433:5
  wire [31:0] _T_3799 = mult_inst198_result + C_reg_bank6_p0_rd_data_2243;	// matmul/matmul-hw.mlir:21225:36, :21420:28, :21434:13
  assign c_i_k_6_i_j_12 = _T_3799;	// matmul/matmul-hw.mlir:21436:5
  //PROBE: c_i_k_6_i_j_12	// matmul/matmul-hw.mlir:21437:5
  assign _T_311 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21438:13
  assign _T_310 = _T_2917 ? _T_3799 : 32'bx;	// matmul/matmul-hw.mlir:8345:18, :21439:13
  localparam [3:0] _T_3801 = 4'h0;	// matmul/matmul-hw.mlir:21442:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21443:5
    if (rst)	// matmul/matmul-hw.mlir:21443:5
      i_k_next_3800 <= _T_3801;	// matmul/matmul-hw.mlir:21446:7
    else	// matmul/matmul-hw.mlir:21443:5
      i_k_next_3800 <= i_k_next_3797;	// matmul/matmul-hw.mlir:21411:13, :21444:7
  end // always @(posedge)
  assign _T_309 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21448:13
  assign _T_308 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21449:13
  mult mult_inst199 (	// matmul/matmul-hw.mlir:21450:28
    .a      (A_reg_bank199_p0_rd_data),	// matmul/matmul-hw.mlir:12414:33
    .b      (_T_2578),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst199_result)
  );
  assign _T_307 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21451:13
  assign a_i_k_7_i_j_12 = A_reg_bank199_p0_rd_data;	// matmul/matmul-hw.mlir:12414:33, :21453:5
  //PROBE: a_i_k_7_i_j_12	// matmul/matmul-hw.mlir:21454:5
  assign b_i_k_7_i_j_12 = _T_2578;	// matmul/matmul-hw.mlir:21456:5
  //PROBE: b_i_k_7_i_j_12	// matmul/matmul-hw.mlir:21457:5
  assign c_prev_i_k_7_i_j_12 = C_reg_bank7_p0_rd_data_2242;	// matmul/matmul-hw.mlir:21226:36, :21459:5
  //PROBE: c_prev_i_k_7_i_j_12	// matmul/matmul-hw.mlir:21460:5
  assign tk_i_k_7_i_j_12 = _T_2902;	// matmul/matmul-hw.mlir:21462:5
  //PROBE: tk_i_k_7_i_j_12	// matmul/matmul-hw.mlir:21463:5
  wire [31:0] _T_3802 = mult_inst199_result + C_reg_bank7_p0_rd_data_2242;	// matmul/matmul-hw.mlir:21226:36, :21450:28, :21464:13
  assign c_i_k_7_i_j_12 = _T_3802;	// matmul/matmul-hw.mlir:21466:5
  //PROBE: c_i_k_7_i_j_12	// matmul/matmul-hw.mlir:21467:5
  assign _T_306 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21468:13
  assign _T_305 = _T_2922 ? _T_3802 : 32'bx;	// matmul/matmul-hw.mlir:8340:18, :21469:13
  localparam [3:0] _T_3804 = 4'h0;	// matmul/matmul-hw.mlir:21472:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21473:5
    if (rst)	// matmul/matmul-hw.mlir:21473:5
      i_k_next_3803 <= _T_3804;	// matmul/matmul-hw.mlir:21476:7
    else	// matmul/matmul-hw.mlir:21473:5
      i_k_next_3803 <= i_k_next_3800;	// matmul/matmul-hw.mlir:21441:13, :21474:7
  end // always @(posedge)
  assign _T_304 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21478:13
  assign _T_303 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21479:13
  mult mult_inst200 (	// matmul/matmul-hw.mlir:21480:28
    .a      (A_reg_bank200_p0_rd_data),	// matmul/matmul-hw.mlir:12415:33
    .b      (_T_2594),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst200_result)
  );
  assign _T_302 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21481:13
  assign a_i_k_8_i_j_12 = A_reg_bank200_p0_rd_data;	// matmul/matmul-hw.mlir:12415:33, :21483:5
  //PROBE: a_i_k_8_i_j_12	// matmul/matmul-hw.mlir:21484:5
  assign b_i_k_8_i_j_12 = _T_2594;	// matmul/matmul-hw.mlir:21486:5
  //PROBE: b_i_k_8_i_j_12	// matmul/matmul-hw.mlir:21487:5
  assign c_prev_i_k_8_i_j_12 = C_reg_bank8_p0_rd_data_2241;	// matmul/matmul-hw.mlir:21227:36, :21489:5
  //PROBE: c_prev_i_k_8_i_j_12	// matmul/matmul-hw.mlir:21490:5
  assign tk_i_k_8_i_j_12 = _T_2907;	// matmul/matmul-hw.mlir:21492:5
  //PROBE: tk_i_k_8_i_j_12	// matmul/matmul-hw.mlir:21493:5
  wire [31:0] _T_3805 = mult_inst200_result + C_reg_bank8_p0_rd_data_2241;	// matmul/matmul-hw.mlir:21227:36, :21480:28, :21494:13
  assign c_i_k_8_i_j_12 = _T_3805;	// matmul/matmul-hw.mlir:21496:5
  //PROBE: c_i_k_8_i_j_12	// matmul/matmul-hw.mlir:21497:5
  assign _T_301 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21498:13
  assign _T_300 = _T_2927 ? _T_3805 : 32'bx;	// matmul/matmul-hw.mlir:8335:18, :21499:13
  localparam [3:0] _T_3807 = 4'h0;	// matmul/matmul-hw.mlir:21502:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21503:5
    if (rst)	// matmul/matmul-hw.mlir:21503:5
      i_k_next_3806 <= _T_3807;	// matmul/matmul-hw.mlir:21506:7
    else	// matmul/matmul-hw.mlir:21503:5
      i_k_next_3806 <= i_k_next_3803;	// matmul/matmul-hw.mlir:21471:13, :21504:7
  end // always @(posedge)
  assign _T_299 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21508:13
  assign _T_298 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21509:13
  mult mult_inst201 (	// matmul/matmul-hw.mlir:21510:28
    .a      (A_reg_bank201_p0_rd_data),	// matmul/matmul-hw.mlir:12416:33
    .b      (_T_2610),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst201_result)
  );
  assign _T_297 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21511:13
  assign a_i_k_9_i_j_12 = A_reg_bank201_p0_rd_data;	// matmul/matmul-hw.mlir:12416:33, :21513:5
  //PROBE: a_i_k_9_i_j_12	// matmul/matmul-hw.mlir:21514:5
  assign b_i_k_9_i_j_12 = _T_2610;	// matmul/matmul-hw.mlir:21516:5
  //PROBE: b_i_k_9_i_j_12	// matmul/matmul-hw.mlir:21517:5
  assign c_prev_i_k_9_i_j_12 = C_reg_bank9_p0_rd_data_2240;	// matmul/matmul-hw.mlir:21228:36, :21519:5
  //PROBE: c_prev_i_k_9_i_j_12	// matmul/matmul-hw.mlir:21520:5
  assign tk_i_k_9_i_j_12 = _T_2912;	// matmul/matmul-hw.mlir:21522:5
  //PROBE: tk_i_k_9_i_j_12	// matmul/matmul-hw.mlir:21523:5
  wire [31:0] _T_3808 = mult_inst201_result + C_reg_bank9_p0_rd_data_2240;	// matmul/matmul-hw.mlir:21228:36, :21510:28, :21524:13
  assign c_i_k_9_i_j_12 = _T_3808;	// matmul/matmul-hw.mlir:21526:5
  //PROBE: c_i_k_9_i_j_12	// matmul/matmul-hw.mlir:21527:5
  assign _T_296 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21528:13
  assign _T_295 = _T_2932 ? _T_3808 : 32'bx;	// matmul/matmul-hw.mlir:8330:18, :21529:13
  localparam [3:0] _T_3810 = 4'h0;	// matmul/matmul-hw.mlir:21532:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21533:5
    if (rst)	// matmul/matmul-hw.mlir:21533:5
      i_k_next_3809 <= _T_3810;	// matmul/matmul-hw.mlir:21536:7
    else	// matmul/matmul-hw.mlir:21533:5
      i_k_next_3809 <= i_k_next_3806;	// matmul/matmul-hw.mlir:21501:13, :21534:7
  end // always @(posedge)
  assign _T_294 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21538:13
  assign _T_293 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21539:13
  mult mult_inst202 (	// matmul/matmul-hw.mlir:21540:28
    .a      (A_reg_bank202_p0_rd_data),	// matmul/matmul-hw.mlir:12417:33
    .b      (_T_2626),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst202_result)
  );
  assign _T_292 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21541:13
  assign a_i_k_10_i_j_12 = A_reg_bank202_p0_rd_data;	// matmul/matmul-hw.mlir:12417:33, :21543:5
  //PROBE: a_i_k_10_i_j_12	// matmul/matmul-hw.mlir:21544:5
  assign b_i_k_10_i_j_12 = _T_2626;	// matmul/matmul-hw.mlir:21546:5
  //PROBE: b_i_k_10_i_j_12	// matmul/matmul-hw.mlir:21547:5
  assign c_prev_i_k_10_i_j_12 = C_reg_bank10_p0_rd_data_2239;	// matmul/matmul-hw.mlir:21229:37, :21549:5
  //PROBE: c_prev_i_k_10_i_j_12	// matmul/matmul-hw.mlir:21550:5
  assign tk_i_k_10_i_j_12 = _T_2917;	// matmul/matmul-hw.mlir:21552:5
  //PROBE: tk_i_k_10_i_j_12	// matmul/matmul-hw.mlir:21553:5
  wire [31:0] _T_3811 = mult_inst202_result + C_reg_bank10_p0_rd_data_2239;	// matmul/matmul-hw.mlir:21229:37, :21540:28, :21554:13
  assign c_i_k_10_i_j_12 = _T_3811;	// matmul/matmul-hw.mlir:21556:5
  //PROBE: c_i_k_10_i_j_12	// matmul/matmul-hw.mlir:21557:5
  assign _T_291 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21558:13
  assign _T_290 = _T_2937 ? _T_3811 : 32'bx;	// matmul/matmul-hw.mlir:8325:18, :21559:13
  localparam [3:0] _T_3813 = 4'h0;	// matmul/matmul-hw.mlir:21562:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21563:5
    if (rst)	// matmul/matmul-hw.mlir:21563:5
      i_k_next_3812 <= _T_3813;	// matmul/matmul-hw.mlir:21566:7
    else	// matmul/matmul-hw.mlir:21563:5
      i_k_next_3812 <= i_k_next_3809;	// matmul/matmul-hw.mlir:21531:13, :21564:7
  end // always @(posedge)
  assign _T_289 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21568:13
  assign _T_288 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21569:13
  mult mult_inst203 (	// matmul/matmul-hw.mlir:21570:28
    .a      (A_reg_bank203_p0_rd_data),	// matmul/matmul-hw.mlir:12418:33
    .b      (_T_2642),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst203_result)
  );
  assign _T_287 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21571:13
  assign a_i_k_11_i_j_12 = A_reg_bank203_p0_rd_data;	// matmul/matmul-hw.mlir:12418:33, :21573:5
  //PROBE: a_i_k_11_i_j_12	// matmul/matmul-hw.mlir:21574:5
  assign b_i_k_11_i_j_12 = _T_2642;	// matmul/matmul-hw.mlir:21576:5
  //PROBE: b_i_k_11_i_j_12	// matmul/matmul-hw.mlir:21577:5
  assign c_prev_i_k_11_i_j_12 = C_reg_bank11_p0_rd_data_2238;	// matmul/matmul-hw.mlir:21230:37, :21579:5
  //PROBE: c_prev_i_k_11_i_j_12	// matmul/matmul-hw.mlir:21580:5
  assign tk_i_k_11_i_j_12 = _T_2922;	// matmul/matmul-hw.mlir:21582:5
  //PROBE: tk_i_k_11_i_j_12	// matmul/matmul-hw.mlir:21583:5
  wire [31:0] _T_3814 = mult_inst203_result + C_reg_bank11_p0_rd_data_2238;	// matmul/matmul-hw.mlir:21230:37, :21570:28, :21584:13
  assign c_i_k_11_i_j_12 = _T_3814;	// matmul/matmul-hw.mlir:21586:5
  //PROBE: c_i_k_11_i_j_12	// matmul/matmul-hw.mlir:21587:5
  assign _T_286 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21588:13
  assign _T_285 = _T_2942 ? _T_3814 : 32'bx;	// matmul/matmul-hw.mlir:8320:18, :21589:13
  localparam [3:0] _T_3816 = 4'h0;	// matmul/matmul-hw.mlir:21592:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21593:5
    if (rst)	// matmul/matmul-hw.mlir:21593:5
      i_k_next_3815 <= _T_3816;	// matmul/matmul-hw.mlir:21596:7
    else	// matmul/matmul-hw.mlir:21593:5
      i_k_next_3815 <= i_k_next_3812;	// matmul/matmul-hw.mlir:21561:13, :21594:7
  end // always @(posedge)
  assign _T_284 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21598:13
  assign _T_283 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21599:13
  mult mult_inst204 (	// matmul/matmul-hw.mlir:21600:28
    .a      (A_reg_bank204_p0_rd_data),	// matmul/matmul-hw.mlir:12419:33
    .b      (_T_2658),
    .t      (_T_2937),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst204_result)
  );
  assign _T_282 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21601:13
  assign a_i_k_12_i_j_12 = A_reg_bank204_p0_rd_data;	// matmul/matmul-hw.mlir:12419:33, :21603:5
  //PROBE: a_i_k_12_i_j_12	// matmul/matmul-hw.mlir:21604:5
  assign b_i_k_12_i_j_12 = _T_2658;	// matmul/matmul-hw.mlir:21606:5
  //PROBE: b_i_k_12_i_j_12	// matmul/matmul-hw.mlir:21607:5
  assign c_prev_i_k_12_i_j_12 = C_reg_bank12_p0_rd_data_2237;	// matmul/matmul-hw.mlir:21231:37, :21609:5
  //PROBE: c_prev_i_k_12_i_j_12	// matmul/matmul-hw.mlir:21610:5
  assign tk_i_k_12_i_j_12 = _T_2927;	// matmul/matmul-hw.mlir:21612:5
  //PROBE: tk_i_k_12_i_j_12	// matmul/matmul-hw.mlir:21613:5
  wire [31:0] _T_3817 = mult_inst204_result + C_reg_bank12_p0_rd_data_2237;	// matmul/matmul-hw.mlir:21231:37, :21600:28, :21614:13
  assign c_i_k_12_i_j_12 = _T_3817;	// matmul/matmul-hw.mlir:21616:5
  //PROBE: c_i_k_12_i_j_12	// matmul/matmul-hw.mlir:21617:5
  assign _T_281 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21618:13
  assign _T_280 = _T_2947 ? _T_3817 : 32'bx;	// matmul/matmul-hw.mlir:8315:18, :21619:13
  localparam [3:0] _T_3819 = 4'h0;	// matmul/matmul-hw.mlir:21622:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21623:5
    if (rst)	// matmul/matmul-hw.mlir:21623:5
      i_k_next_3818 <= _T_3819;	// matmul/matmul-hw.mlir:21626:7
    else	// matmul/matmul-hw.mlir:21623:5
      i_k_next_3818 <= i_k_next_3815;	// matmul/matmul-hw.mlir:21591:13, :21624:7
  end // always @(posedge)
  assign _T_279 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21628:13
  assign _T_278 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21629:13
  mult mult_inst205 (	// matmul/matmul-hw.mlir:21630:28
    .a      (A_reg_bank205_p0_rd_data),	// matmul/matmul-hw.mlir:12420:33
    .b      (_T_2674),
    .t      (_T_2942),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst205_result)
  );
  assign _T_277 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21631:13
  assign a_i_k_13_i_j_12 = A_reg_bank205_p0_rd_data;	// matmul/matmul-hw.mlir:12420:33, :21633:5
  //PROBE: a_i_k_13_i_j_12	// matmul/matmul-hw.mlir:21634:5
  assign b_i_k_13_i_j_12 = _T_2674;	// matmul/matmul-hw.mlir:21636:5
  //PROBE: b_i_k_13_i_j_12	// matmul/matmul-hw.mlir:21637:5
  assign c_prev_i_k_13_i_j_12 = C_reg_bank13_p0_rd_data_2236;	// matmul/matmul-hw.mlir:21232:37, :21639:5
  //PROBE: c_prev_i_k_13_i_j_12	// matmul/matmul-hw.mlir:21640:5
  assign tk_i_k_13_i_j_12 = _T_2932;	// matmul/matmul-hw.mlir:21642:5
  //PROBE: tk_i_k_13_i_j_12	// matmul/matmul-hw.mlir:21643:5
  wire [31:0] _T_3820 = mult_inst205_result + C_reg_bank13_p0_rd_data_2236;	// matmul/matmul-hw.mlir:21232:37, :21630:28, :21644:13
  assign c_i_k_13_i_j_12 = _T_3820;	// matmul/matmul-hw.mlir:21646:5
  //PROBE: c_i_k_13_i_j_12	// matmul/matmul-hw.mlir:21647:5
  assign _T_276 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21648:13
  assign _T_275 = _T_2952 ? _T_3820 : 32'bx;	// matmul/matmul-hw.mlir:8310:18, :21649:13
  localparam [3:0] _T_3822 = 4'h0;	// matmul/matmul-hw.mlir:21652:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21653:5
    if (rst)	// matmul/matmul-hw.mlir:21653:5
      i_k_next_3821 <= _T_3822;	// matmul/matmul-hw.mlir:21656:7
    else	// matmul/matmul-hw.mlir:21653:5
      i_k_next_3821 <= i_k_next_3818;	// matmul/matmul-hw.mlir:21621:13, :21654:7
  end // always @(posedge)
  assign _T_274 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21658:13
  assign _T_273 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21659:13
  mult mult_inst206 (	// matmul/matmul-hw.mlir:21660:28
    .a      (A_reg_bank206_p0_rd_data),	// matmul/matmul-hw.mlir:12421:33
    .b      (_T_2690),
    .t      (_T_2947),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst206_result)
  );
  assign _T_272 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21661:13
  assign a_i_k_14_i_j_12 = A_reg_bank206_p0_rd_data;	// matmul/matmul-hw.mlir:12421:33, :21663:5
  //PROBE: a_i_k_14_i_j_12	// matmul/matmul-hw.mlir:21664:5
  assign b_i_k_14_i_j_12 = _T_2690;	// matmul/matmul-hw.mlir:21666:5
  //PROBE: b_i_k_14_i_j_12	// matmul/matmul-hw.mlir:21667:5
  assign c_prev_i_k_14_i_j_12 = C_reg_bank14_p0_rd_data_2235;	// matmul/matmul-hw.mlir:21233:37, :21669:5
  //PROBE: c_prev_i_k_14_i_j_12	// matmul/matmul-hw.mlir:21670:5
  assign tk_i_k_14_i_j_12 = _T_2937;	// matmul/matmul-hw.mlir:21672:5
  //PROBE: tk_i_k_14_i_j_12	// matmul/matmul-hw.mlir:21673:5
  wire [31:0] _T_3823 = mult_inst206_result + C_reg_bank14_p0_rd_data_2235;	// matmul/matmul-hw.mlir:21233:37, :21660:28, :21674:13
  assign c_i_k_14_i_j_12 = _T_3823;	// matmul/matmul-hw.mlir:21676:5
  //PROBE: c_i_k_14_i_j_12	// matmul/matmul-hw.mlir:21677:5
  assign _T_271 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21678:13
  assign _T_270 = _T_2957 ? _T_3823 : 32'bx;	// matmul/matmul-hw.mlir:8305:18, :21679:13
  localparam [3:0] _T_3825 = 4'h0;	// matmul/matmul-hw.mlir:21682:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21683:5
    if (rst)	// matmul/matmul-hw.mlir:21683:5
      i_k_next_3824 <= _T_3825;	// matmul/matmul-hw.mlir:21686:7
    else	// matmul/matmul-hw.mlir:21683:5
      i_k_next_3824 <= i_k_next_3821;	// matmul/matmul-hw.mlir:21651:13, :21684:7
  end // always @(posedge)
  assign _T_269 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21688:13
  assign _T_268 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21689:13
  mult mult_inst207 (	// matmul/matmul-hw.mlir:21690:28
    .a      (A_reg_bank207_p0_rd_data),	// matmul/matmul-hw.mlir:12422:33
    .b      (_T_2706),
    .t      (_T_2952),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst207_result)
  );
  assign _T_267 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21691:13
  assign a_i_k_15_i_j_12 = A_reg_bank207_p0_rd_data;	// matmul/matmul-hw.mlir:12422:33, :21693:5
  //PROBE: a_i_k_15_i_j_12	// matmul/matmul-hw.mlir:21694:5
  assign b_i_k_15_i_j_12 = _T_2706;	// matmul/matmul-hw.mlir:21696:5
  //PROBE: b_i_k_15_i_j_12	// matmul/matmul-hw.mlir:21697:5
  assign c_prev_i_k_15_i_j_12 = C_reg_bank15_p0_rd_data_2234;	// matmul/matmul-hw.mlir:21234:37, :21699:5
  //PROBE: c_prev_i_k_15_i_j_12	// matmul/matmul-hw.mlir:21700:5
  assign tk_i_k_15_i_j_12 = _T_2942;	// matmul/matmul-hw.mlir:21702:5
  //PROBE: tk_i_k_15_i_j_12	// matmul/matmul-hw.mlir:21703:5
  wire [31:0] _T_3826 = mult_inst207_result + C_reg_bank15_p0_rd_data_2234;	// matmul/matmul-hw.mlir:21234:37, :21690:28, :21704:13
  assign c_i_k_15_i_j_12 = _T_3826;	// matmul/matmul-hw.mlir:21706:5
  //PROBE: c_i_k_15_i_j_12	// matmul/matmul-hw.mlir:21707:5
  assign _T_266 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21708:13
  assign _T_265 = _T_2962 ? _T_3826 : 32'bx;	// matmul/matmul-hw.mlir:8300:18, :21709:13
  localparam [3:0] _T_3828 = 4'h0;	// matmul/matmul-hw.mlir:21712:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21713:5
    if (rst)	// matmul/matmul-hw.mlir:21713:5
      i_k_next_3827 <= _T_3828;	// matmul/matmul-hw.mlir:21716:7
    else	// matmul/matmul-hw.mlir:21713:5
      i_k_next_3827 <= i_k_next_3824;	// matmul/matmul-hw.mlir:21681:13, :21714:7
  end // always @(posedge)
  wire [31:0] _T_3830 = _T_3829;	// matmul/matmul-hw.mlir:21719:13
  wire [31:0] _T_3831 = {_T_3830[5'h0+:31], {{_T_2712}}};	// matmul/matmul-hw.mlir:21720:19, :21721:13, :21722:13, :21723:13
  wire [31:0] _T_3832 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:21724:19, :21725:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21726:5
    if (rst)	// matmul/matmul-hw.mlir:21726:5
      _T_3829 <= _T_3832;	// matmul/matmul-hw.mlir:21729:7
    else	// matmul/matmul-hw.mlir:21726:5
      _T_3829 <= _T_3831;	// matmul/matmul-hw.mlir:21727:7
  end // always @(posedge)
  wire _T_3833 = _T_3829[5'h1F];	// matmul/matmul-hw.mlir:21719:13, :21731:15, :21732:13
  assign _T_264 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21733:13
  wire [3:0][3:0] _T_3835 = i_delayed_3834;	// matmul/matmul-hw.mlir:21735:13
  wire [3:0][3:0] _T_3836 = {_T_3835[2'h0+:3], {{i_k_next_3827}}};	// matmul/matmul-hw.mlir:21711:13, :21736:19, :21737:13, :21738:13, :21739:13
  wire [3:0][3:0] _T_3837 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:21740:19, :21741:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21742:5
    if (rst)	// matmul/matmul-hw.mlir:21742:5
      i_delayed_3834 <= _T_3837;	// matmul/matmul-hw.mlir:21745:7
    else	// matmul/matmul-hw.mlir:21742:5
      i_delayed_3834 <= _T_3836;	// matmul/matmul-hw.mlir:21743:7
  end // always @(posedge)
  assign _T_263 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21749:13
  assign _T_262 = _T_3833 ? i_delayed_3834[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8297:17, :21735:13, :21747:20, :21748:13, :21750:13
  assign _T_261 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21751:13
  assign _T_260 = _T_3833 ? C_reg_bank16_p0_rd_data_2233 : 32'bx;	// matmul/matmul-hw.mlir:8295:18, :21235:37, :21752:13
  localparam [3:0] _T_3839 = 4'h0;	// matmul/matmul-hw.mlir:21755:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21756:5
    if (rst)	// matmul/matmul-hw.mlir:21756:5
      i_j_next_3838 <= _T_3839;	// matmul/matmul-hw.mlir:21759:7
    else	// matmul/matmul-hw.mlir:21756:5
      i_j_next_3838 <= i_j_next_3762;	// matmul/matmul-hw.mlir:21144:13, :21757:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3840 (	// matmul/matmul-hw.mlir:21829:36
    .p0_rd_en   (_T_255),	// matmul/matmul-hw.mlir:21851:13
    .p1_wr_en   (_T_259),	// matmul/matmul-hw.mlir:21846:13
    .p1_wr_data (_T_258),	// matmul/matmul-hw.mlir:21847:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2232)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3841 (	// matmul/matmul-hw.mlir:21830:36
    .p0_rd_en   (_T_250),	// matmul/matmul-hw.mlir:21881:13
    .p1_wr_en   (_T_254),	// matmul/matmul-hw.mlir:21868:13
    .p1_wr_data (_T_253),	// matmul/matmul-hw.mlir:21869:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2231)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3842 (	// matmul/matmul-hw.mlir:21831:36
    .p0_rd_en   (_T_245),	// matmul/matmul-hw.mlir:21911:13
    .p1_wr_en   (_T_249),	// matmul/matmul-hw.mlir:21898:13
    .p1_wr_data (_T_248),	// matmul/matmul-hw.mlir:21899:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2230)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3843 (	// matmul/matmul-hw.mlir:21832:36
    .p0_rd_en   (_T_240),	// matmul/matmul-hw.mlir:21941:13
    .p1_wr_en   (_T_244),	// matmul/matmul-hw.mlir:21928:13
    .p1_wr_data (_T_243),	// matmul/matmul-hw.mlir:21929:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2229)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3844 (	// matmul/matmul-hw.mlir:21833:36
    .p0_rd_en   (_T_235),	// matmul/matmul-hw.mlir:21971:13
    .p1_wr_en   (_T_239),	// matmul/matmul-hw.mlir:21958:13
    .p1_wr_data (_T_238),	// matmul/matmul-hw.mlir:21959:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2228)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3845 (	// matmul/matmul-hw.mlir:21834:36
    .p0_rd_en   (_T_230),	// matmul/matmul-hw.mlir:22001:13
    .p1_wr_en   (_T_234),	// matmul/matmul-hw.mlir:21988:13
    .p1_wr_data (_T_233),	// matmul/matmul-hw.mlir:21989:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2227)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3846 (	// matmul/matmul-hw.mlir:21835:36
    .p0_rd_en   (_T_225),	// matmul/matmul-hw.mlir:22031:13
    .p1_wr_en   (_T_229),	// matmul/matmul-hw.mlir:22018:13
    .p1_wr_data (_T_228),	// matmul/matmul-hw.mlir:22019:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2226)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3847 (	// matmul/matmul-hw.mlir:21836:36
    .p0_rd_en   (_T_220),	// matmul/matmul-hw.mlir:22061:13
    .p1_wr_en   (_T_224),	// matmul/matmul-hw.mlir:22048:13
    .p1_wr_data (_T_223),	// matmul/matmul-hw.mlir:22049:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2225)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3848 (	// matmul/matmul-hw.mlir:21837:36
    .p0_rd_en   (_T_215),	// matmul/matmul-hw.mlir:22091:13
    .p1_wr_en   (_T_219),	// matmul/matmul-hw.mlir:22078:13
    .p1_wr_data (_T_218),	// matmul/matmul-hw.mlir:22079:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2224)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3849 (	// matmul/matmul-hw.mlir:21838:36
    .p0_rd_en   (_T_210),	// matmul/matmul-hw.mlir:22121:13
    .p1_wr_en   (_T_214),	// matmul/matmul-hw.mlir:22108:13
    .p1_wr_data (_T_213),	// matmul/matmul-hw.mlir:22109:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2223)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3850 (	// matmul/matmul-hw.mlir:21839:37
    .p0_rd_en   (_T_205),	// matmul/matmul-hw.mlir:22151:13
    .p1_wr_en   (_T_209),	// matmul/matmul-hw.mlir:22138:13
    .p1_wr_data (_T_208),	// matmul/matmul-hw.mlir:22139:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2222)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3851 (	// matmul/matmul-hw.mlir:21840:37
    .p0_rd_en   (_T_200),	// matmul/matmul-hw.mlir:22181:13
    .p1_wr_en   (_T_204),	// matmul/matmul-hw.mlir:22168:13
    .p1_wr_data (_T_203),	// matmul/matmul-hw.mlir:22169:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2221)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3852 (	// matmul/matmul-hw.mlir:21841:37
    .p0_rd_en   (_T_195),	// matmul/matmul-hw.mlir:22211:13
    .p1_wr_en   (_T_199),	// matmul/matmul-hw.mlir:22198:13
    .p1_wr_data (_T_198),	// matmul/matmul-hw.mlir:22199:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2220)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3853 (	// matmul/matmul-hw.mlir:21842:37
    .p0_rd_en   (_T_190),	// matmul/matmul-hw.mlir:22241:13
    .p1_wr_en   (_T_194),	// matmul/matmul-hw.mlir:22228:13
    .p1_wr_data (_T_193),	// matmul/matmul-hw.mlir:22229:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2219)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3854 (	// matmul/matmul-hw.mlir:21843:37
    .p0_rd_en   (_T_185),	// matmul/matmul-hw.mlir:22271:13
    .p1_wr_en   (_T_189),	// matmul/matmul-hw.mlir:22258:13
    .p1_wr_data (_T_188),	// matmul/matmul-hw.mlir:22259:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2218)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3855 (	// matmul/matmul-hw.mlir:21844:37
    .p0_rd_en   (_T_180),	// matmul/matmul-hw.mlir:22301:13
    .p1_wr_en   (_T_184),	// matmul/matmul-hw.mlir:22288:13
    .p1_wr_data (_T_183),	// matmul/matmul-hw.mlir:22289:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2217)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3856 (	// matmul/matmul-hw.mlir:21845:37
    .p0_rd_en   (_T_177),	// matmul/matmul-hw.mlir:22343:13
    .p1_wr_en   (_T_179),	// matmul/matmul-hw.mlir:22318:13
    .p1_wr_data (_T_178),	// matmul/matmul-hw.mlir:22319:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2216)
  );
  assign _T_259 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21846:13
  assign _T_258 = _T_2885 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8293:18, :21847:13
  assign _T_257 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21848:13
  assign _T_256 = _T_2874 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21849:13
  mult mult_inst208 (	// matmul/matmul-hw.mlir:21850:28
    .a      (A_reg_bank208_p0_rd_data),	// matmul/matmul-hw.mlir:12423:33
    .b      (_T_2467),
    .t      (_T_2874),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst208_result)
  );
  assign _T_255 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21851:13
  assign a_i_k_0_i_j_13 = A_reg_bank208_p0_rd_data;	// matmul/matmul-hw.mlir:12423:33, :21853:5
  //PROBE: a_i_k_0_i_j_13	// matmul/matmul-hw.mlir:21854:5
  assign b_i_k_0_i_j_13 = _T_2467;	// matmul/matmul-hw.mlir:21856:5
  //PROBE: b_i_k_0_i_j_13	// matmul/matmul-hw.mlir:21857:5
  assign c_prev_i_k_0_i_j_13 = C_reg_bank0_p0_rd_data_2232;	// matmul/matmul-hw.mlir:21829:36, :21859:5
  //PROBE: c_prev_i_k_0_i_j_13	// matmul/matmul-hw.mlir:21860:5
  assign tk_i_k_0_i_j_13 = _T_2852;	// matmul/matmul-hw.mlir:21862:5
  //PROBE: tk_i_k_0_i_j_13	// matmul/matmul-hw.mlir:21863:5
  wire [31:0] _T_3857 = mult_inst208_result + C_reg_bank0_p0_rd_data_2232;	// matmul/matmul-hw.mlir:21829:36, :21850:28, :21864:13
  assign c_i_k_0_i_j_13 = _T_3857;	// matmul/matmul-hw.mlir:21866:5
  //PROBE: c_i_k_0_i_j_13	// matmul/matmul-hw.mlir:21867:5
  assign _T_254 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21868:13
  assign _T_253 = _T_2892 ? _T_3857 : 32'bx;	// matmul/matmul-hw.mlir:8288:18, :21869:13
  localparam [3:0] _T_3859 = 4'h0;	// matmul/matmul-hw.mlir:21872:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21873:5
    if (rst)	// matmul/matmul-hw.mlir:21873:5
      i_k_next_3858 <= _T_3859;	// matmul/matmul-hw.mlir:21876:7
    else	// matmul/matmul-hw.mlir:21873:5
      i_k_next_3858 <= i_j_next_3838;	// matmul/matmul-hw.mlir:21754:13, :21874:7
  end // always @(posedge)
  assign _T_252 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21878:13
  assign _T_251 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21879:13
  mult mult_inst209 (	// matmul/matmul-hw.mlir:21880:28
    .a      (A_reg_bank209_p0_rd_data),	// matmul/matmul-hw.mlir:12424:33
    .b      (_T_2483),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst209_result)
  );
  assign _T_250 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21881:13
  assign a_i_k_1_i_j_13 = A_reg_bank209_p0_rd_data;	// matmul/matmul-hw.mlir:12424:33, :21883:5
  //PROBE: a_i_k_1_i_j_13	// matmul/matmul-hw.mlir:21884:5
  assign b_i_k_1_i_j_13 = _T_2483;	// matmul/matmul-hw.mlir:21886:5
  //PROBE: b_i_k_1_i_j_13	// matmul/matmul-hw.mlir:21887:5
  assign c_prev_i_k_1_i_j_13 = C_reg_bank1_p0_rd_data_2231;	// matmul/matmul-hw.mlir:21830:36, :21889:5
  //PROBE: c_prev_i_k_1_i_j_13	// matmul/matmul-hw.mlir:21890:5
  assign tk_i_k_1_i_j_13 = _T_2863;	// matmul/matmul-hw.mlir:21892:5
  //PROBE: tk_i_k_1_i_j_13	// matmul/matmul-hw.mlir:21893:5
  wire [31:0] _T_3860 = mult_inst209_result + C_reg_bank1_p0_rd_data_2231;	// matmul/matmul-hw.mlir:21830:36, :21880:28, :21894:13
  assign c_i_k_1_i_j_13 = _T_3860;	// matmul/matmul-hw.mlir:21896:5
  //PROBE: c_i_k_1_i_j_13	// matmul/matmul-hw.mlir:21897:5
  assign _T_249 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21898:13
  assign _T_248 = _T_2897 ? _T_3860 : 32'bx;	// matmul/matmul-hw.mlir:8283:18, :21899:13
  localparam [3:0] _T_3862 = 4'h0;	// matmul/matmul-hw.mlir:21902:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21903:5
    if (rst)	// matmul/matmul-hw.mlir:21903:5
      i_k_next_3861 <= _T_3862;	// matmul/matmul-hw.mlir:21906:7
    else	// matmul/matmul-hw.mlir:21903:5
      i_k_next_3861 <= i_k_next_3858;	// matmul/matmul-hw.mlir:21871:13, :21904:7
  end // always @(posedge)
  assign _T_247 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21908:13
  assign _T_246 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21909:13
  mult mult_inst210 (	// matmul/matmul-hw.mlir:21910:28
    .a      (A_reg_bank210_p0_rd_data),	// matmul/matmul-hw.mlir:12425:33
    .b      (_T_2499),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst210_result)
  );
  assign _T_245 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21911:13
  assign a_i_k_2_i_j_13 = A_reg_bank210_p0_rd_data;	// matmul/matmul-hw.mlir:12425:33, :21913:5
  //PROBE: a_i_k_2_i_j_13	// matmul/matmul-hw.mlir:21914:5
  assign b_i_k_2_i_j_13 = _T_2499;	// matmul/matmul-hw.mlir:21916:5
  //PROBE: b_i_k_2_i_j_13	// matmul/matmul-hw.mlir:21917:5
  assign c_prev_i_k_2_i_j_13 = C_reg_bank2_p0_rd_data_2230;	// matmul/matmul-hw.mlir:21831:36, :21919:5
  //PROBE: c_prev_i_k_2_i_j_13	// matmul/matmul-hw.mlir:21920:5
  assign tk_i_k_2_i_j_13 = _T_2874;	// matmul/matmul-hw.mlir:21922:5
  //PROBE: tk_i_k_2_i_j_13	// matmul/matmul-hw.mlir:21923:5
  wire [31:0] _T_3863 = mult_inst210_result + C_reg_bank2_p0_rd_data_2230;	// matmul/matmul-hw.mlir:21831:36, :21910:28, :21924:13
  assign c_i_k_2_i_j_13 = _T_3863;	// matmul/matmul-hw.mlir:21926:5
  //PROBE: c_i_k_2_i_j_13	// matmul/matmul-hw.mlir:21927:5
  assign _T_244 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21928:13
  assign _T_243 = _T_2902 ? _T_3863 : 32'bx;	// matmul/matmul-hw.mlir:8278:18, :21929:13
  localparam [3:0] _T_3865 = 4'h0;	// matmul/matmul-hw.mlir:21932:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21933:5
    if (rst)	// matmul/matmul-hw.mlir:21933:5
      i_k_next_3864 <= _T_3865;	// matmul/matmul-hw.mlir:21936:7
    else	// matmul/matmul-hw.mlir:21933:5
      i_k_next_3864 <= i_k_next_3861;	// matmul/matmul-hw.mlir:21901:13, :21934:7
  end // always @(posedge)
  assign _T_242 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21938:13
  assign _T_241 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21939:13
  mult mult_inst211 (	// matmul/matmul-hw.mlir:21940:28
    .a      (A_reg_bank211_p0_rd_data),	// matmul/matmul-hw.mlir:12426:33
    .b      (_T_2515),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst211_result)
  );
  assign _T_240 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21941:13
  assign a_i_k_3_i_j_13 = A_reg_bank211_p0_rd_data;	// matmul/matmul-hw.mlir:12426:33, :21943:5
  //PROBE: a_i_k_3_i_j_13	// matmul/matmul-hw.mlir:21944:5
  assign b_i_k_3_i_j_13 = _T_2515;	// matmul/matmul-hw.mlir:21946:5
  //PROBE: b_i_k_3_i_j_13	// matmul/matmul-hw.mlir:21947:5
  assign c_prev_i_k_3_i_j_13 = C_reg_bank3_p0_rd_data_2229;	// matmul/matmul-hw.mlir:21832:36, :21949:5
  //PROBE: c_prev_i_k_3_i_j_13	// matmul/matmul-hw.mlir:21950:5
  assign tk_i_k_3_i_j_13 = _T_2885;	// matmul/matmul-hw.mlir:21952:5
  //PROBE: tk_i_k_3_i_j_13	// matmul/matmul-hw.mlir:21953:5
  wire [31:0] _T_3866 = mult_inst211_result + C_reg_bank3_p0_rd_data_2229;	// matmul/matmul-hw.mlir:21832:36, :21940:28, :21954:13
  assign c_i_k_3_i_j_13 = _T_3866;	// matmul/matmul-hw.mlir:21956:5
  //PROBE: c_i_k_3_i_j_13	// matmul/matmul-hw.mlir:21957:5
  assign _T_239 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21958:13
  assign _T_238 = _T_2907 ? _T_3866 : 32'bx;	// matmul/matmul-hw.mlir:8273:18, :21959:13
  localparam [3:0] _T_3868 = 4'h0;	// matmul/matmul-hw.mlir:21962:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21963:5
    if (rst)	// matmul/matmul-hw.mlir:21963:5
      i_k_next_3867 <= _T_3868;	// matmul/matmul-hw.mlir:21966:7
    else	// matmul/matmul-hw.mlir:21963:5
      i_k_next_3867 <= i_k_next_3864;	// matmul/matmul-hw.mlir:21931:13, :21964:7
  end // always @(posedge)
  assign _T_237 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21968:13
  assign _T_236 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21969:13
  mult mult_inst212 (	// matmul/matmul-hw.mlir:21970:28
    .a      (A_reg_bank212_p0_rd_data),	// matmul/matmul-hw.mlir:12427:33
    .b      (_T_2531),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst212_result)
  );
  assign _T_235 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21971:13
  assign a_i_k_4_i_j_13 = A_reg_bank212_p0_rd_data;	// matmul/matmul-hw.mlir:12427:33, :21973:5
  //PROBE: a_i_k_4_i_j_13	// matmul/matmul-hw.mlir:21974:5
  assign b_i_k_4_i_j_13 = _T_2531;	// matmul/matmul-hw.mlir:21976:5
  //PROBE: b_i_k_4_i_j_13	// matmul/matmul-hw.mlir:21977:5
  assign c_prev_i_k_4_i_j_13 = C_reg_bank4_p0_rd_data_2228;	// matmul/matmul-hw.mlir:21833:36, :21979:5
  //PROBE: c_prev_i_k_4_i_j_13	// matmul/matmul-hw.mlir:21980:5
  assign tk_i_k_4_i_j_13 = _T_2892;	// matmul/matmul-hw.mlir:21982:5
  //PROBE: tk_i_k_4_i_j_13	// matmul/matmul-hw.mlir:21983:5
  wire [31:0] _T_3869 = mult_inst212_result + C_reg_bank4_p0_rd_data_2228;	// matmul/matmul-hw.mlir:21833:36, :21970:28, :21984:13
  assign c_i_k_4_i_j_13 = _T_3869;	// matmul/matmul-hw.mlir:21986:5
  //PROBE: c_i_k_4_i_j_13	// matmul/matmul-hw.mlir:21987:5
  assign _T_234 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21988:13
  assign _T_233 = _T_2912 ? _T_3869 : 32'bx;	// matmul/matmul-hw.mlir:8268:18, :21989:13
  localparam [3:0] _T_3871 = 4'h0;	// matmul/matmul-hw.mlir:21992:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:21993:5
    if (rst)	// matmul/matmul-hw.mlir:21993:5
      i_k_next_3870 <= _T_3871;	// matmul/matmul-hw.mlir:21996:7
    else	// matmul/matmul-hw.mlir:21993:5
      i_k_next_3870 <= i_k_next_3867;	// matmul/matmul-hw.mlir:21961:13, :21994:7
  end // always @(posedge)
  assign _T_232 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21998:13
  assign _T_231 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :21999:13
  mult mult_inst213 (	// matmul/matmul-hw.mlir:22000:28
    .a      (A_reg_bank213_p0_rd_data),	// matmul/matmul-hw.mlir:12428:33
    .b      (_T_2547),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst213_result)
  );
  assign _T_230 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22001:13
  assign a_i_k_5_i_j_13 = A_reg_bank213_p0_rd_data;	// matmul/matmul-hw.mlir:12428:33, :22003:5
  //PROBE: a_i_k_5_i_j_13	// matmul/matmul-hw.mlir:22004:5
  assign b_i_k_5_i_j_13 = _T_2547;	// matmul/matmul-hw.mlir:22006:5
  //PROBE: b_i_k_5_i_j_13	// matmul/matmul-hw.mlir:22007:5
  assign c_prev_i_k_5_i_j_13 = C_reg_bank5_p0_rd_data_2227;	// matmul/matmul-hw.mlir:21834:36, :22009:5
  //PROBE: c_prev_i_k_5_i_j_13	// matmul/matmul-hw.mlir:22010:5
  assign tk_i_k_5_i_j_13 = _T_2897;	// matmul/matmul-hw.mlir:22012:5
  //PROBE: tk_i_k_5_i_j_13	// matmul/matmul-hw.mlir:22013:5
  wire [31:0] _T_3872 = mult_inst213_result + C_reg_bank5_p0_rd_data_2227;	// matmul/matmul-hw.mlir:21834:36, :22000:28, :22014:13
  assign c_i_k_5_i_j_13 = _T_3872;	// matmul/matmul-hw.mlir:22016:5
  //PROBE: c_i_k_5_i_j_13	// matmul/matmul-hw.mlir:22017:5
  assign _T_229 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22018:13
  assign _T_228 = _T_2917 ? _T_3872 : 32'bx;	// matmul/matmul-hw.mlir:8263:18, :22019:13
  localparam [3:0] _T_3874 = 4'h0;	// matmul/matmul-hw.mlir:22022:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22023:5
    if (rst)	// matmul/matmul-hw.mlir:22023:5
      i_k_next_3873 <= _T_3874;	// matmul/matmul-hw.mlir:22026:7
    else	// matmul/matmul-hw.mlir:22023:5
      i_k_next_3873 <= i_k_next_3870;	// matmul/matmul-hw.mlir:21991:13, :22024:7
  end // always @(posedge)
  assign _T_227 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22028:13
  assign _T_226 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22029:13
  mult mult_inst214 (	// matmul/matmul-hw.mlir:22030:28
    .a      (A_reg_bank214_p0_rd_data),	// matmul/matmul-hw.mlir:12429:33
    .b      (_T_2563),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst214_result)
  );
  assign _T_225 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22031:13
  assign a_i_k_6_i_j_13 = A_reg_bank214_p0_rd_data;	// matmul/matmul-hw.mlir:12429:33, :22033:5
  //PROBE: a_i_k_6_i_j_13	// matmul/matmul-hw.mlir:22034:5
  assign b_i_k_6_i_j_13 = _T_2563;	// matmul/matmul-hw.mlir:22036:5
  //PROBE: b_i_k_6_i_j_13	// matmul/matmul-hw.mlir:22037:5
  assign c_prev_i_k_6_i_j_13 = C_reg_bank6_p0_rd_data_2226;	// matmul/matmul-hw.mlir:21835:36, :22039:5
  //PROBE: c_prev_i_k_6_i_j_13	// matmul/matmul-hw.mlir:22040:5
  assign tk_i_k_6_i_j_13 = _T_2902;	// matmul/matmul-hw.mlir:22042:5
  //PROBE: tk_i_k_6_i_j_13	// matmul/matmul-hw.mlir:22043:5
  wire [31:0] _T_3875 = mult_inst214_result + C_reg_bank6_p0_rd_data_2226;	// matmul/matmul-hw.mlir:21835:36, :22030:28, :22044:13
  assign c_i_k_6_i_j_13 = _T_3875;	// matmul/matmul-hw.mlir:22046:5
  //PROBE: c_i_k_6_i_j_13	// matmul/matmul-hw.mlir:22047:5
  assign _T_224 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22048:13
  assign _T_223 = _T_2922 ? _T_3875 : 32'bx;	// matmul/matmul-hw.mlir:8258:18, :22049:13
  localparam [3:0] _T_3877 = 4'h0;	// matmul/matmul-hw.mlir:22052:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22053:5
    if (rst)	// matmul/matmul-hw.mlir:22053:5
      i_k_next_3876 <= _T_3877;	// matmul/matmul-hw.mlir:22056:7
    else	// matmul/matmul-hw.mlir:22053:5
      i_k_next_3876 <= i_k_next_3873;	// matmul/matmul-hw.mlir:22021:13, :22054:7
  end // always @(posedge)
  assign _T_222 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22058:13
  assign _T_221 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22059:13
  mult mult_inst215 (	// matmul/matmul-hw.mlir:22060:28
    .a      (A_reg_bank215_p0_rd_data),	// matmul/matmul-hw.mlir:12430:33
    .b      (_T_2579),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst215_result)
  );
  assign _T_220 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22061:13
  assign a_i_k_7_i_j_13 = A_reg_bank215_p0_rd_data;	// matmul/matmul-hw.mlir:12430:33, :22063:5
  //PROBE: a_i_k_7_i_j_13	// matmul/matmul-hw.mlir:22064:5
  assign b_i_k_7_i_j_13 = _T_2579;	// matmul/matmul-hw.mlir:22066:5
  //PROBE: b_i_k_7_i_j_13	// matmul/matmul-hw.mlir:22067:5
  assign c_prev_i_k_7_i_j_13 = C_reg_bank7_p0_rd_data_2225;	// matmul/matmul-hw.mlir:21836:36, :22069:5
  //PROBE: c_prev_i_k_7_i_j_13	// matmul/matmul-hw.mlir:22070:5
  assign tk_i_k_7_i_j_13 = _T_2907;	// matmul/matmul-hw.mlir:22072:5
  //PROBE: tk_i_k_7_i_j_13	// matmul/matmul-hw.mlir:22073:5
  wire [31:0] _T_3878 = mult_inst215_result + C_reg_bank7_p0_rd_data_2225;	// matmul/matmul-hw.mlir:21836:36, :22060:28, :22074:13
  assign c_i_k_7_i_j_13 = _T_3878;	// matmul/matmul-hw.mlir:22076:5
  //PROBE: c_i_k_7_i_j_13	// matmul/matmul-hw.mlir:22077:5
  assign _T_219 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22078:13
  assign _T_218 = _T_2927 ? _T_3878 : 32'bx;	// matmul/matmul-hw.mlir:8253:18, :22079:13
  localparam [3:0] _T_3880 = 4'h0;	// matmul/matmul-hw.mlir:22082:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22083:5
    if (rst)	// matmul/matmul-hw.mlir:22083:5
      i_k_next_3879 <= _T_3880;	// matmul/matmul-hw.mlir:22086:7
    else	// matmul/matmul-hw.mlir:22083:5
      i_k_next_3879 <= i_k_next_3876;	// matmul/matmul-hw.mlir:22051:13, :22084:7
  end // always @(posedge)
  assign _T_217 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22088:13
  assign _T_216 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22089:13
  mult mult_inst216 (	// matmul/matmul-hw.mlir:22090:28
    .a      (A_reg_bank216_p0_rd_data),	// matmul/matmul-hw.mlir:12431:33
    .b      (_T_2595),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst216_result)
  );
  assign _T_215 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22091:13
  assign a_i_k_8_i_j_13 = A_reg_bank216_p0_rd_data;	// matmul/matmul-hw.mlir:12431:33, :22093:5
  //PROBE: a_i_k_8_i_j_13	// matmul/matmul-hw.mlir:22094:5
  assign b_i_k_8_i_j_13 = _T_2595;	// matmul/matmul-hw.mlir:22096:5
  //PROBE: b_i_k_8_i_j_13	// matmul/matmul-hw.mlir:22097:5
  assign c_prev_i_k_8_i_j_13 = C_reg_bank8_p0_rd_data_2224;	// matmul/matmul-hw.mlir:21837:36, :22099:5
  //PROBE: c_prev_i_k_8_i_j_13	// matmul/matmul-hw.mlir:22100:5
  assign tk_i_k_8_i_j_13 = _T_2912;	// matmul/matmul-hw.mlir:22102:5
  //PROBE: tk_i_k_8_i_j_13	// matmul/matmul-hw.mlir:22103:5
  wire [31:0] _T_3881 = mult_inst216_result + C_reg_bank8_p0_rd_data_2224;	// matmul/matmul-hw.mlir:21837:36, :22090:28, :22104:13
  assign c_i_k_8_i_j_13 = _T_3881;	// matmul/matmul-hw.mlir:22106:5
  //PROBE: c_i_k_8_i_j_13	// matmul/matmul-hw.mlir:22107:5
  assign _T_214 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22108:13
  assign _T_213 = _T_2932 ? _T_3881 : 32'bx;	// matmul/matmul-hw.mlir:8248:18, :22109:13
  localparam [3:0] _T_3883 = 4'h0;	// matmul/matmul-hw.mlir:22112:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22113:5
    if (rst)	// matmul/matmul-hw.mlir:22113:5
      i_k_next_3882 <= _T_3883;	// matmul/matmul-hw.mlir:22116:7
    else	// matmul/matmul-hw.mlir:22113:5
      i_k_next_3882 <= i_k_next_3879;	// matmul/matmul-hw.mlir:22081:13, :22114:7
  end // always @(posedge)
  assign _T_212 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22118:13
  assign _T_211 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22119:13
  mult mult_inst217 (	// matmul/matmul-hw.mlir:22120:28
    .a      (A_reg_bank217_p0_rd_data),	// matmul/matmul-hw.mlir:12432:33
    .b      (_T_2611),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst217_result)
  );
  assign _T_210 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22121:13
  assign a_i_k_9_i_j_13 = A_reg_bank217_p0_rd_data;	// matmul/matmul-hw.mlir:12432:33, :22123:5
  //PROBE: a_i_k_9_i_j_13	// matmul/matmul-hw.mlir:22124:5
  assign b_i_k_9_i_j_13 = _T_2611;	// matmul/matmul-hw.mlir:22126:5
  //PROBE: b_i_k_9_i_j_13	// matmul/matmul-hw.mlir:22127:5
  assign c_prev_i_k_9_i_j_13 = C_reg_bank9_p0_rd_data_2223;	// matmul/matmul-hw.mlir:21838:36, :22129:5
  //PROBE: c_prev_i_k_9_i_j_13	// matmul/matmul-hw.mlir:22130:5
  assign tk_i_k_9_i_j_13 = _T_2917;	// matmul/matmul-hw.mlir:22132:5
  //PROBE: tk_i_k_9_i_j_13	// matmul/matmul-hw.mlir:22133:5
  wire [31:0] _T_3884 = mult_inst217_result + C_reg_bank9_p0_rd_data_2223;	// matmul/matmul-hw.mlir:21838:36, :22120:28, :22134:13
  assign c_i_k_9_i_j_13 = _T_3884;	// matmul/matmul-hw.mlir:22136:5
  //PROBE: c_i_k_9_i_j_13	// matmul/matmul-hw.mlir:22137:5
  assign _T_209 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22138:13
  assign _T_208 = _T_2937 ? _T_3884 : 32'bx;	// matmul/matmul-hw.mlir:8243:18, :22139:13
  localparam [3:0] _T_3886 = 4'h0;	// matmul/matmul-hw.mlir:22142:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22143:5
    if (rst)	// matmul/matmul-hw.mlir:22143:5
      i_k_next_3885 <= _T_3886;	// matmul/matmul-hw.mlir:22146:7
    else	// matmul/matmul-hw.mlir:22143:5
      i_k_next_3885 <= i_k_next_3882;	// matmul/matmul-hw.mlir:22111:13, :22144:7
  end // always @(posedge)
  assign _T_207 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22148:13
  assign _T_206 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22149:13
  mult mult_inst218 (	// matmul/matmul-hw.mlir:22150:28
    .a      (A_reg_bank218_p0_rd_data),	// matmul/matmul-hw.mlir:12433:33
    .b      (_T_2627),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst218_result)
  );
  assign _T_205 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22151:13
  assign a_i_k_10_i_j_13 = A_reg_bank218_p0_rd_data;	// matmul/matmul-hw.mlir:12433:33, :22153:5
  //PROBE: a_i_k_10_i_j_13	// matmul/matmul-hw.mlir:22154:5
  assign b_i_k_10_i_j_13 = _T_2627;	// matmul/matmul-hw.mlir:22156:5
  //PROBE: b_i_k_10_i_j_13	// matmul/matmul-hw.mlir:22157:5
  assign c_prev_i_k_10_i_j_13 = C_reg_bank10_p0_rd_data_2222;	// matmul/matmul-hw.mlir:21839:37, :22159:5
  //PROBE: c_prev_i_k_10_i_j_13	// matmul/matmul-hw.mlir:22160:5
  assign tk_i_k_10_i_j_13 = _T_2922;	// matmul/matmul-hw.mlir:22162:5
  //PROBE: tk_i_k_10_i_j_13	// matmul/matmul-hw.mlir:22163:5
  wire [31:0] _T_3887 = mult_inst218_result + C_reg_bank10_p0_rd_data_2222;	// matmul/matmul-hw.mlir:21839:37, :22150:28, :22164:13
  assign c_i_k_10_i_j_13 = _T_3887;	// matmul/matmul-hw.mlir:22166:5
  //PROBE: c_i_k_10_i_j_13	// matmul/matmul-hw.mlir:22167:5
  assign _T_204 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22168:13
  assign _T_203 = _T_2942 ? _T_3887 : 32'bx;	// matmul/matmul-hw.mlir:8238:18, :22169:13
  localparam [3:0] _T_3889 = 4'h0;	// matmul/matmul-hw.mlir:22172:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22173:5
    if (rst)	// matmul/matmul-hw.mlir:22173:5
      i_k_next_3888 <= _T_3889;	// matmul/matmul-hw.mlir:22176:7
    else	// matmul/matmul-hw.mlir:22173:5
      i_k_next_3888 <= i_k_next_3885;	// matmul/matmul-hw.mlir:22141:13, :22174:7
  end // always @(posedge)
  assign _T_202 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22178:13
  assign _T_201 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22179:13
  mult mult_inst219 (	// matmul/matmul-hw.mlir:22180:28
    .a      (A_reg_bank219_p0_rd_data),	// matmul/matmul-hw.mlir:12434:33
    .b      (_T_2643),
    .t      (_T_2937),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst219_result)
  );
  assign _T_200 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22181:13
  assign a_i_k_11_i_j_13 = A_reg_bank219_p0_rd_data;	// matmul/matmul-hw.mlir:12434:33, :22183:5
  //PROBE: a_i_k_11_i_j_13	// matmul/matmul-hw.mlir:22184:5
  assign b_i_k_11_i_j_13 = _T_2643;	// matmul/matmul-hw.mlir:22186:5
  //PROBE: b_i_k_11_i_j_13	// matmul/matmul-hw.mlir:22187:5
  assign c_prev_i_k_11_i_j_13 = C_reg_bank11_p0_rd_data_2221;	// matmul/matmul-hw.mlir:21840:37, :22189:5
  //PROBE: c_prev_i_k_11_i_j_13	// matmul/matmul-hw.mlir:22190:5
  assign tk_i_k_11_i_j_13 = _T_2927;	// matmul/matmul-hw.mlir:22192:5
  //PROBE: tk_i_k_11_i_j_13	// matmul/matmul-hw.mlir:22193:5
  wire [31:0] _T_3890 = mult_inst219_result + C_reg_bank11_p0_rd_data_2221;	// matmul/matmul-hw.mlir:21840:37, :22180:28, :22194:13
  assign c_i_k_11_i_j_13 = _T_3890;	// matmul/matmul-hw.mlir:22196:5
  //PROBE: c_i_k_11_i_j_13	// matmul/matmul-hw.mlir:22197:5
  assign _T_199 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22198:13
  assign _T_198 = _T_2947 ? _T_3890 : 32'bx;	// matmul/matmul-hw.mlir:8233:18, :22199:13
  localparam [3:0] _T_3892 = 4'h0;	// matmul/matmul-hw.mlir:22202:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22203:5
    if (rst)	// matmul/matmul-hw.mlir:22203:5
      i_k_next_3891 <= _T_3892;	// matmul/matmul-hw.mlir:22206:7
    else	// matmul/matmul-hw.mlir:22203:5
      i_k_next_3891 <= i_k_next_3888;	// matmul/matmul-hw.mlir:22171:13, :22204:7
  end // always @(posedge)
  assign _T_197 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22208:13
  assign _T_196 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22209:13
  mult mult_inst220 (	// matmul/matmul-hw.mlir:22210:28
    .a      (A_reg_bank220_p0_rd_data),	// matmul/matmul-hw.mlir:12435:33
    .b      (_T_2659),
    .t      (_T_2942),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst220_result)
  );
  assign _T_195 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22211:13
  assign a_i_k_12_i_j_13 = A_reg_bank220_p0_rd_data;	// matmul/matmul-hw.mlir:12435:33, :22213:5
  //PROBE: a_i_k_12_i_j_13	// matmul/matmul-hw.mlir:22214:5
  assign b_i_k_12_i_j_13 = _T_2659;	// matmul/matmul-hw.mlir:22216:5
  //PROBE: b_i_k_12_i_j_13	// matmul/matmul-hw.mlir:22217:5
  assign c_prev_i_k_12_i_j_13 = C_reg_bank12_p0_rd_data_2220;	// matmul/matmul-hw.mlir:21841:37, :22219:5
  //PROBE: c_prev_i_k_12_i_j_13	// matmul/matmul-hw.mlir:22220:5
  assign tk_i_k_12_i_j_13 = _T_2932;	// matmul/matmul-hw.mlir:22222:5
  //PROBE: tk_i_k_12_i_j_13	// matmul/matmul-hw.mlir:22223:5
  wire [31:0] _T_3893 = mult_inst220_result + C_reg_bank12_p0_rd_data_2220;	// matmul/matmul-hw.mlir:21841:37, :22210:28, :22224:13
  assign c_i_k_12_i_j_13 = _T_3893;	// matmul/matmul-hw.mlir:22226:5
  //PROBE: c_i_k_12_i_j_13	// matmul/matmul-hw.mlir:22227:5
  assign _T_194 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22228:13
  assign _T_193 = _T_2952 ? _T_3893 : 32'bx;	// matmul/matmul-hw.mlir:8228:18, :22229:13
  localparam [3:0] _T_3895 = 4'h0;	// matmul/matmul-hw.mlir:22232:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22233:5
    if (rst)	// matmul/matmul-hw.mlir:22233:5
      i_k_next_3894 <= _T_3895;	// matmul/matmul-hw.mlir:22236:7
    else	// matmul/matmul-hw.mlir:22233:5
      i_k_next_3894 <= i_k_next_3891;	// matmul/matmul-hw.mlir:22201:13, :22234:7
  end // always @(posedge)
  assign _T_192 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22238:13
  assign _T_191 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22239:13
  mult mult_inst221 (	// matmul/matmul-hw.mlir:22240:28
    .a      (A_reg_bank221_p0_rd_data),	// matmul/matmul-hw.mlir:12436:33
    .b      (_T_2675),
    .t      (_T_2947),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst221_result)
  );
  assign _T_190 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22241:13
  assign a_i_k_13_i_j_13 = A_reg_bank221_p0_rd_data;	// matmul/matmul-hw.mlir:12436:33, :22243:5
  //PROBE: a_i_k_13_i_j_13	// matmul/matmul-hw.mlir:22244:5
  assign b_i_k_13_i_j_13 = _T_2675;	// matmul/matmul-hw.mlir:22246:5
  //PROBE: b_i_k_13_i_j_13	// matmul/matmul-hw.mlir:22247:5
  assign c_prev_i_k_13_i_j_13 = C_reg_bank13_p0_rd_data_2219;	// matmul/matmul-hw.mlir:21842:37, :22249:5
  //PROBE: c_prev_i_k_13_i_j_13	// matmul/matmul-hw.mlir:22250:5
  assign tk_i_k_13_i_j_13 = _T_2937;	// matmul/matmul-hw.mlir:22252:5
  //PROBE: tk_i_k_13_i_j_13	// matmul/matmul-hw.mlir:22253:5
  wire [31:0] _T_3896 = mult_inst221_result + C_reg_bank13_p0_rd_data_2219;	// matmul/matmul-hw.mlir:21842:37, :22240:28, :22254:13
  assign c_i_k_13_i_j_13 = _T_3896;	// matmul/matmul-hw.mlir:22256:5
  //PROBE: c_i_k_13_i_j_13	// matmul/matmul-hw.mlir:22257:5
  assign _T_189 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22258:13
  assign _T_188 = _T_2957 ? _T_3896 : 32'bx;	// matmul/matmul-hw.mlir:8223:18, :22259:13
  localparam [3:0] _T_3898 = 4'h0;	// matmul/matmul-hw.mlir:22262:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22263:5
    if (rst)	// matmul/matmul-hw.mlir:22263:5
      i_k_next_3897 <= _T_3898;	// matmul/matmul-hw.mlir:22266:7
    else	// matmul/matmul-hw.mlir:22263:5
      i_k_next_3897 <= i_k_next_3894;	// matmul/matmul-hw.mlir:22231:13, :22264:7
  end // always @(posedge)
  assign _T_187 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22268:13
  assign _T_186 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22269:13
  mult mult_inst222 (	// matmul/matmul-hw.mlir:22270:28
    .a      (A_reg_bank222_p0_rd_data),	// matmul/matmul-hw.mlir:12437:33
    .b      (_T_2691),
    .t      (_T_2952),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst222_result)
  );
  assign _T_185 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22271:13
  assign a_i_k_14_i_j_13 = A_reg_bank222_p0_rd_data;	// matmul/matmul-hw.mlir:12437:33, :22273:5
  //PROBE: a_i_k_14_i_j_13	// matmul/matmul-hw.mlir:22274:5
  assign b_i_k_14_i_j_13 = _T_2691;	// matmul/matmul-hw.mlir:22276:5
  //PROBE: b_i_k_14_i_j_13	// matmul/matmul-hw.mlir:22277:5
  assign c_prev_i_k_14_i_j_13 = C_reg_bank14_p0_rd_data_2218;	// matmul/matmul-hw.mlir:21843:37, :22279:5
  //PROBE: c_prev_i_k_14_i_j_13	// matmul/matmul-hw.mlir:22280:5
  assign tk_i_k_14_i_j_13 = _T_2942;	// matmul/matmul-hw.mlir:22282:5
  //PROBE: tk_i_k_14_i_j_13	// matmul/matmul-hw.mlir:22283:5
  wire [31:0] _T_3899 = mult_inst222_result + C_reg_bank14_p0_rd_data_2218;	// matmul/matmul-hw.mlir:21843:37, :22270:28, :22284:13
  assign c_i_k_14_i_j_13 = _T_3899;	// matmul/matmul-hw.mlir:22286:5
  //PROBE: c_i_k_14_i_j_13	// matmul/matmul-hw.mlir:22287:5
  assign _T_184 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22288:13
  assign _T_183 = _T_2962 ? _T_3899 : 32'bx;	// matmul/matmul-hw.mlir:8218:18, :22289:13
  localparam [3:0] _T_3901 = 4'h0;	// matmul/matmul-hw.mlir:22292:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22293:5
    if (rst)	// matmul/matmul-hw.mlir:22293:5
      i_k_next_3900 <= _T_3901;	// matmul/matmul-hw.mlir:22296:7
    else	// matmul/matmul-hw.mlir:22293:5
      i_k_next_3900 <= i_k_next_3897;	// matmul/matmul-hw.mlir:22261:13, :22294:7
  end // always @(posedge)
  assign _T_182 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22298:13
  assign _T_181 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22299:13
  mult mult_inst223 (	// matmul/matmul-hw.mlir:22300:28
    .a      (A_reg_bank223_p0_rd_data),	// matmul/matmul-hw.mlir:12438:33
    .b      (_T_2707),
    .t      (_T_2957),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst223_result)
  );
  assign _T_180 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22301:13
  assign a_i_k_15_i_j_13 = A_reg_bank223_p0_rd_data;	// matmul/matmul-hw.mlir:12438:33, :22303:5
  //PROBE: a_i_k_15_i_j_13	// matmul/matmul-hw.mlir:22304:5
  assign b_i_k_15_i_j_13 = _T_2707;	// matmul/matmul-hw.mlir:22306:5
  //PROBE: b_i_k_15_i_j_13	// matmul/matmul-hw.mlir:22307:5
  assign c_prev_i_k_15_i_j_13 = C_reg_bank15_p0_rd_data_2217;	// matmul/matmul-hw.mlir:21844:37, :22309:5
  //PROBE: c_prev_i_k_15_i_j_13	// matmul/matmul-hw.mlir:22310:5
  assign tk_i_k_15_i_j_13 = _T_2947;	// matmul/matmul-hw.mlir:22312:5
  //PROBE: tk_i_k_15_i_j_13	// matmul/matmul-hw.mlir:22313:5
  wire [31:0] _T_3902 = mult_inst223_result + C_reg_bank15_p0_rd_data_2217;	// matmul/matmul-hw.mlir:21844:37, :22300:28, :22314:13
  assign c_i_k_15_i_j_13 = _T_3902;	// matmul/matmul-hw.mlir:22316:5
  //PROBE: c_i_k_15_i_j_13	// matmul/matmul-hw.mlir:22317:5
  assign _T_179 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22318:13
  assign _T_178 = _T_3833 ? _T_3902 : 32'bx;	// matmul/matmul-hw.mlir:8213:18, :22319:13
  localparam [3:0] _T_3904 = 4'h0;	// matmul/matmul-hw.mlir:22322:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22323:5
    if (rst)	// matmul/matmul-hw.mlir:22323:5
      i_k_next_3903 <= _T_3904;	// matmul/matmul-hw.mlir:22326:7
    else	// matmul/matmul-hw.mlir:22323:5
      i_k_next_3903 <= i_k_next_3900;	// matmul/matmul-hw.mlir:22291:13, :22324:7
  end // always @(posedge)
  wire [32:0] _T_3906 = _T_3905;	// matmul/matmul-hw.mlir:22329:13
  wire [32:0] _T_3907 = {_T_3906[6'h0+:32], {{_T_2712}}};	// matmul/matmul-hw.mlir:22330:19, :22331:13, :22332:13, :22333:13
  wire [32:0] _T_3908 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:22334:19, :22335:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22336:5
    if (rst)	// matmul/matmul-hw.mlir:22336:5
      _T_3905 <= _T_3908;	// matmul/matmul-hw.mlir:22339:7
    else	// matmul/matmul-hw.mlir:22336:5
      _T_3905 <= _T_3907;	// matmul/matmul-hw.mlir:22337:7
  end // always @(posedge)
  wire _T_3909 = _T_3905[6'h20];	// matmul/matmul-hw.mlir:22329:13, :22341:16, :22342:13
  assign _T_177 = _T_3909 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22343:13
  wire [3:0][3:0] _T_3911 = i_delayed_3910;	// matmul/matmul-hw.mlir:22345:13
  wire [3:0][3:0] _T_3912 = {_T_3911[2'h0+:3], {{i_k_next_3903}}};	// matmul/matmul-hw.mlir:22321:13, :22346:19, :22347:13, :22348:13, :22349:13
  wire [3:0][3:0] _T_3913 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:22350:19, :22351:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22352:5
    if (rst)	// matmul/matmul-hw.mlir:22352:5
      i_delayed_3910 <= _T_3913;	// matmul/matmul-hw.mlir:22355:7
    else	// matmul/matmul-hw.mlir:22352:5
      i_delayed_3910 <= _T_3912;	// matmul/matmul-hw.mlir:22353:7
  end // always @(posedge)
  assign _T_176 = _T_3909 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22359:13
  assign _T_175 = _T_3909 ? i_delayed_3910[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8210:17, :22345:13, :22357:20, :22358:13, :22360:13
  assign _T_174 = _T_3909 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22361:13
  assign _T_173 = _T_3909 ? C_reg_bank16_p0_rd_data_2216 : 32'bx;	// matmul/matmul-hw.mlir:8208:18, :21845:37, :22362:13
  localparam [3:0] _T_3915 = 4'h0;	// matmul/matmul-hw.mlir:22365:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22366:5
    if (rst)	// matmul/matmul-hw.mlir:22366:5
      i_j_next_3914 <= _T_3915;	// matmul/matmul-hw.mlir:22369:7
    else	// matmul/matmul-hw.mlir:22366:5
      i_j_next_3914 <= i_j_next_3838;	// matmul/matmul-hw.mlir:21754:13, :22367:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3916 (	// matmul/matmul-hw.mlir:22439:36
    .p0_rd_en   (_T_168),	// matmul/matmul-hw.mlir:22461:13
    .p1_wr_en   (_T_172),	// matmul/matmul-hw.mlir:22456:13
    .p1_wr_data (_T_171),	// matmul/matmul-hw.mlir:22457:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data_2215)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3917 (	// matmul/matmul-hw.mlir:22440:36
    .p0_rd_en   (_T_163),	// matmul/matmul-hw.mlir:22491:13
    .p1_wr_en   (_T_167),	// matmul/matmul-hw.mlir:22478:13
    .p1_wr_data (_T_166),	// matmul/matmul-hw.mlir:22479:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data_2214)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3918 (	// matmul/matmul-hw.mlir:22441:36
    .p0_rd_en   (_T_158),	// matmul/matmul-hw.mlir:22521:13
    .p1_wr_en   (_T_162),	// matmul/matmul-hw.mlir:22508:13
    .p1_wr_data (_T_161),	// matmul/matmul-hw.mlir:22509:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data_2213)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3919 (	// matmul/matmul-hw.mlir:22442:36
    .p0_rd_en   (_T_153),	// matmul/matmul-hw.mlir:22551:13
    .p1_wr_en   (_T_157),	// matmul/matmul-hw.mlir:22538:13
    .p1_wr_data (_T_156),	// matmul/matmul-hw.mlir:22539:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data_2212)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3920 (	// matmul/matmul-hw.mlir:22443:36
    .p0_rd_en   (_T_148),	// matmul/matmul-hw.mlir:22581:13
    .p1_wr_en   (_T_152),	// matmul/matmul-hw.mlir:22568:13
    .p1_wr_data (_T_151),	// matmul/matmul-hw.mlir:22569:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data_2211)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3921 (	// matmul/matmul-hw.mlir:22444:36
    .p0_rd_en   (_T_143),	// matmul/matmul-hw.mlir:22611:13
    .p1_wr_en   (_T_147),	// matmul/matmul-hw.mlir:22598:13
    .p1_wr_data (_T_146),	// matmul/matmul-hw.mlir:22599:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data_2210)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3922 (	// matmul/matmul-hw.mlir:22445:36
    .p0_rd_en   (_T_138),	// matmul/matmul-hw.mlir:22641:13
    .p1_wr_en   (_T_142),	// matmul/matmul-hw.mlir:22628:13
    .p1_wr_data (_T_141),	// matmul/matmul-hw.mlir:22629:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data_2209)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3923 (	// matmul/matmul-hw.mlir:22446:36
    .p0_rd_en   (_T_133),	// matmul/matmul-hw.mlir:22671:13
    .p1_wr_en   (_T_137),	// matmul/matmul-hw.mlir:22658:13
    .p1_wr_data (_T_136),	// matmul/matmul-hw.mlir:22659:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data_2208)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_3924 (	// matmul/matmul-hw.mlir:22447:36
    .p0_rd_en   (_T_128),	// matmul/matmul-hw.mlir:22701:13
    .p1_wr_en   (_T_132),	// matmul/matmul-hw.mlir:22688:13
    .p1_wr_data (_T_131),	// matmul/matmul-hw.mlir:22689:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data_2207)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_3925 (	// matmul/matmul-hw.mlir:22448:36
    .p0_rd_en   (_T_123),	// matmul/matmul-hw.mlir:22731:13
    .p1_wr_en   (_T_127),	// matmul/matmul-hw.mlir:22718:13
    .p1_wr_data (_T_126),	// matmul/matmul-hw.mlir:22719:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data_2206)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_3926 (	// matmul/matmul-hw.mlir:22449:37
    .p0_rd_en   (_T_118),	// matmul/matmul-hw.mlir:22761:13
    .p1_wr_en   (_T_122),	// matmul/matmul-hw.mlir:22748:13
    .p1_wr_data (_T_121),	// matmul/matmul-hw.mlir:22749:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data_2205)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_3927 (	// matmul/matmul-hw.mlir:22450:37
    .p0_rd_en   (_T_113),	// matmul/matmul-hw.mlir:22791:13
    .p1_wr_en   (_T_117),	// matmul/matmul-hw.mlir:22778:13
    .p1_wr_data (_T_116),	// matmul/matmul-hw.mlir:22779:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data_2204)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_3928 (	// matmul/matmul-hw.mlir:22451:37
    .p0_rd_en   (_T_108),	// matmul/matmul-hw.mlir:22821:13
    .p1_wr_en   (_T_112),	// matmul/matmul-hw.mlir:22808:13
    .p1_wr_data (_T_111),	// matmul/matmul-hw.mlir:22809:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data_2203)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_3929 (	// matmul/matmul-hw.mlir:22452:37
    .p0_rd_en   (_T_103),	// matmul/matmul-hw.mlir:22851:13
    .p1_wr_en   (_T_107),	// matmul/matmul-hw.mlir:22838:13
    .p1_wr_data (_T_106),	// matmul/matmul-hw.mlir:22839:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data_2202)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_3930 (	// matmul/matmul-hw.mlir:22453:37
    .p0_rd_en   (_T_98),	// matmul/matmul-hw.mlir:22881:13
    .p1_wr_en   (_T_102),	// matmul/matmul-hw.mlir:22868:13
    .p1_wr_data (_T_101),	// matmul/matmul-hw.mlir:22869:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data_2201)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_3931 (	// matmul/matmul-hw.mlir:22454:37
    .p0_rd_en   (_T_93),	// matmul/matmul-hw.mlir:22911:13
    .p1_wr_en   (_T_97),	// matmul/matmul-hw.mlir:22898:13
    .p1_wr_data (_T_96),	// matmul/matmul-hw.mlir:22899:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data_2200)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_3932 (	// matmul/matmul-hw.mlir:22455:37
    .p0_rd_en   (_T_90),	// matmul/matmul-hw.mlir:22953:13
    .p1_wr_en   (_T_92),	// matmul/matmul-hw.mlir:22928:13
    .p1_wr_data (_T_91),	// matmul/matmul-hw.mlir:22929:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data_2199)
  );
  assign _T_172 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22456:13
  assign _T_171 = _T_2892 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8206:18, :22457:13
  assign _T_170 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22458:13
  assign _T_169 = _T_2885 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22459:13
  mult mult_inst224 (	// matmul/matmul-hw.mlir:22460:28
    .a      (A_reg_bank224_p0_rd_data),	// matmul/matmul-hw.mlir:12439:33
    .b      (_T_2468),
    .t      (_T_2885),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst224_result)
  );
  assign _T_168 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22461:13
  assign a_i_k_0_i_j_14 = A_reg_bank224_p0_rd_data;	// matmul/matmul-hw.mlir:12439:33, :22463:5
  //PROBE: a_i_k_0_i_j_14	// matmul/matmul-hw.mlir:22464:5
  assign b_i_k_0_i_j_14 = _T_2468;	// matmul/matmul-hw.mlir:22466:5
  //PROBE: b_i_k_0_i_j_14	// matmul/matmul-hw.mlir:22467:5
  assign c_prev_i_k_0_i_j_14 = C_reg_bank0_p0_rd_data_2215;	// matmul/matmul-hw.mlir:22439:36, :22469:5
  //PROBE: c_prev_i_k_0_i_j_14	// matmul/matmul-hw.mlir:22470:5
  assign tk_i_k_0_i_j_14 = _T_2863;	// matmul/matmul-hw.mlir:22472:5
  //PROBE: tk_i_k_0_i_j_14	// matmul/matmul-hw.mlir:22473:5
  wire [31:0] _T_3933 = mult_inst224_result + C_reg_bank0_p0_rd_data_2215;	// matmul/matmul-hw.mlir:22439:36, :22460:28, :22474:13
  assign c_i_k_0_i_j_14 = _T_3933;	// matmul/matmul-hw.mlir:22476:5
  //PROBE: c_i_k_0_i_j_14	// matmul/matmul-hw.mlir:22477:5
  assign _T_167 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22478:13
  assign _T_166 = _T_2897 ? _T_3933 : 32'bx;	// matmul/matmul-hw.mlir:8201:18, :22479:13
  localparam [3:0] _T_3935 = 4'h0;	// matmul/matmul-hw.mlir:22482:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22483:5
    if (rst)	// matmul/matmul-hw.mlir:22483:5
      i_k_next_3934 <= _T_3935;	// matmul/matmul-hw.mlir:22486:7
    else	// matmul/matmul-hw.mlir:22483:5
      i_k_next_3934 <= i_j_next_3914;	// matmul/matmul-hw.mlir:22364:13, :22484:7
  end // always @(posedge)
  assign _T_165 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22488:13
  assign _T_164 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22489:13
  mult mult_inst225 (	// matmul/matmul-hw.mlir:22490:28
    .a      (A_reg_bank225_p0_rd_data),	// matmul/matmul-hw.mlir:12440:33
    .b      (_T_2484),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst225_result)
  );
  assign _T_163 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22491:13
  assign a_i_k_1_i_j_14 = A_reg_bank225_p0_rd_data;	// matmul/matmul-hw.mlir:12440:33, :22493:5
  //PROBE: a_i_k_1_i_j_14	// matmul/matmul-hw.mlir:22494:5
  assign b_i_k_1_i_j_14 = _T_2484;	// matmul/matmul-hw.mlir:22496:5
  //PROBE: b_i_k_1_i_j_14	// matmul/matmul-hw.mlir:22497:5
  assign c_prev_i_k_1_i_j_14 = C_reg_bank1_p0_rd_data_2214;	// matmul/matmul-hw.mlir:22440:36, :22499:5
  //PROBE: c_prev_i_k_1_i_j_14	// matmul/matmul-hw.mlir:22500:5
  assign tk_i_k_1_i_j_14 = _T_2874;	// matmul/matmul-hw.mlir:22502:5
  //PROBE: tk_i_k_1_i_j_14	// matmul/matmul-hw.mlir:22503:5
  wire [31:0] _T_3936 = mult_inst225_result + C_reg_bank1_p0_rd_data_2214;	// matmul/matmul-hw.mlir:22440:36, :22490:28, :22504:13
  assign c_i_k_1_i_j_14 = _T_3936;	// matmul/matmul-hw.mlir:22506:5
  //PROBE: c_i_k_1_i_j_14	// matmul/matmul-hw.mlir:22507:5
  assign _T_162 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22508:13
  assign _T_161 = _T_2902 ? _T_3936 : 32'bx;	// matmul/matmul-hw.mlir:8196:18, :22509:13
  localparam [3:0] _T_3938 = 4'h0;	// matmul/matmul-hw.mlir:22512:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22513:5
    if (rst)	// matmul/matmul-hw.mlir:22513:5
      i_k_next_3937 <= _T_3938;	// matmul/matmul-hw.mlir:22516:7
    else	// matmul/matmul-hw.mlir:22513:5
      i_k_next_3937 <= i_k_next_3934;	// matmul/matmul-hw.mlir:22481:13, :22514:7
  end // always @(posedge)
  assign _T_160 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22518:13
  assign _T_159 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22519:13
  mult mult_inst226 (	// matmul/matmul-hw.mlir:22520:28
    .a      (A_reg_bank226_p0_rd_data),	// matmul/matmul-hw.mlir:12441:33
    .b      (_T_2500),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst226_result)
  );
  assign _T_158 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22521:13
  assign a_i_k_2_i_j_14 = A_reg_bank226_p0_rd_data;	// matmul/matmul-hw.mlir:12441:33, :22523:5
  //PROBE: a_i_k_2_i_j_14	// matmul/matmul-hw.mlir:22524:5
  assign b_i_k_2_i_j_14 = _T_2500;	// matmul/matmul-hw.mlir:22526:5
  //PROBE: b_i_k_2_i_j_14	// matmul/matmul-hw.mlir:22527:5
  assign c_prev_i_k_2_i_j_14 = C_reg_bank2_p0_rd_data_2213;	// matmul/matmul-hw.mlir:22441:36, :22529:5
  //PROBE: c_prev_i_k_2_i_j_14	// matmul/matmul-hw.mlir:22530:5
  assign tk_i_k_2_i_j_14 = _T_2885;	// matmul/matmul-hw.mlir:22532:5
  //PROBE: tk_i_k_2_i_j_14	// matmul/matmul-hw.mlir:22533:5
  wire [31:0] _T_3939 = mult_inst226_result + C_reg_bank2_p0_rd_data_2213;	// matmul/matmul-hw.mlir:22441:36, :22520:28, :22534:13
  assign c_i_k_2_i_j_14 = _T_3939;	// matmul/matmul-hw.mlir:22536:5
  //PROBE: c_i_k_2_i_j_14	// matmul/matmul-hw.mlir:22537:5
  assign _T_157 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22538:13
  assign _T_156 = _T_2907 ? _T_3939 : 32'bx;	// matmul/matmul-hw.mlir:8191:18, :22539:13
  localparam [3:0] _T_3941 = 4'h0;	// matmul/matmul-hw.mlir:22542:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22543:5
    if (rst)	// matmul/matmul-hw.mlir:22543:5
      i_k_next_3940 <= _T_3941;	// matmul/matmul-hw.mlir:22546:7
    else	// matmul/matmul-hw.mlir:22543:5
      i_k_next_3940 <= i_k_next_3937;	// matmul/matmul-hw.mlir:22511:13, :22544:7
  end // always @(posedge)
  assign _T_155 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22548:13
  assign _T_154 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22549:13
  mult mult_inst227 (	// matmul/matmul-hw.mlir:22550:28
    .a      (A_reg_bank227_p0_rd_data),	// matmul/matmul-hw.mlir:12442:33
    .b      (_T_2516),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst227_result)
  );
  assign _T_153 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22551:13
  assign a_i_k_3_i_j_14 = A_reg_bank227_p0_rd_data;	// matmul/matmul-hw.mlir:12442:33, :22553:5
  //PROBE: a_i_k_3_i_j_14	// matmul/matmul-hw.mlir:22554:5
  assign b_i_k_3_i_j_14 = _T_2516;	// matmul/matmul-hw.mlir:22556:5
  //PROBE: b_i_k_3_i_j_14	// matmul/matmul-hw.mlir:22557:5
  assign c_prev_i_k_3_i_j_14 = C_reg_bank3_p0_rd_data_2212;	// matmul/matmul-hw.mlir:22442:36, :22559:5
  //PROBE: c_prev_i_k_3_i_j_14	// matmul/matmul-hw.mlir:22560:5
  assign tk_i_k_3_i_j_14 = _T_2892;	// matmul/matmul-hw.mlir:22562:5
  //PROBE: tk_i_k_3_i_j_14	// matmul/matmul-hw.mlir:22563:5
  wire [31:0] _T_3942 = mult_inst227_result + C_reg_bank3_p0_rd_data_2212;	// matmul/matmul-hw.mlir:22442:36, :22550:28, :22564:13
  assign c_i_k_3_i_j_14 = _T_3942;	// matmul/matmul-hw.mlir:22566:5
  //PROBE: c_i_k_3_i_j_14	// matmul/matmul-hw.mlir:22567:5
  assign _T_152 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22568:13
  assign _T_151 = _T_2912 ? _T_3942 : 32'bx;	// matmul/matmul-hw.mlir:8186:18, :22569:13
  localparam [3:0] _T_3944 = 4'h0;	// matmul/matmul-hw.mlir:22572:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22573:5
    if (rst)	// matmul/matmul-hw.mlir:22573:5
      i_k_next_3943 <= _T_3944;	// matmul/matmul-hw.mlir:22576:7
    else	// matmul/matmul-hw.mlir:22573:5
      i_k_next_3943 <= i_k_next_3940;	// matmul/matmul-hw.mlir:22541:13, :22574:7
  end // always @(posedge)
  assign _T_150 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22578:13
  assign _T_149 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22579:13
  mult mult_inst228 (	// matmul/matmul-hw.mlir:22580:28
    .a      (A_reg_bank228_p0_rd_data),	// matmul/matmul-hw.mlir:12443:33
    .b      (_T_2532),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst228_result)
  );
  assign _T_148 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22581:13
  assign a_i_k_4_i_j_14 = A_reg_bank228_p0_rd_data;	// matmul/matmul-hw.mlir:12443:33, :22583:5
  //PROBE: a_i_k_4_i_j_14	// matmul/matmul-hw.mlir:22584:5
  assign b_i_k_4_i_j_14 = _T_2532;	// matmul/matmul-hw.mlir:22586:5
  //PROBE: b_i_k_4_i_j_14	// matmul/matmul-hw.mlir:22587:5
  assign c_prev_i_k_4_i_j_14 = C_reg_bank4_p0_rd_data_2211;	// matmul/matmul-hw.mlir:22443:36, :22589:5
  //PROBE: c_prev_i_k_4_i_j_14	// matmul/matmul-hw.mlir:22590:5
  assign tk_i_k_4_i_j_14 = _T_2897;	// matmul/matmul-hw.mlir:22592:5
  //PROBE: tk_i_k_4_i_j_14	// matmul/matmul-hw.mlir:22593:5
  wire [31:0] _T_3945 = mult_inst228_result + C_reg_bank4_p0_rd_data_2211;	// matmul/matmul-hw.mlir:22443:36, :22580:28, :22594:13
  assign c_i_k_4_i_j_14 = _T_3945;	// matmul/matmul-hw.mlir:22596:5
  //PROBE: c_i_k_4_i_j_14	// matmul/matmul-hw.mlir:22597:5
  assign _T_147 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22598:13
  assign _T_146 = _T_2917 ? _T_3945 : 32'bx;	// matmul/matmul-hw.mlir:8181:18, :22599:13
  localparam [3:0] _T_3947 = 4'h0;	// matmul/matmul-hw.mlir:22602:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22603:5
    if (rst)	// matmul/matmul-hw.mlir:22603:5
      i_k_next_3946 <= _T_3947;	// matmul/matmul-hw.mlir:22606:7
    else	// matmul/matmul-hw.mlir:22603:5
      i_k_next_3946 <= i_k_next_3943;	// matmul/matmul-hw.mlir:22571:13, :22604:7
  end // always @(posedge)
  assign _T_145 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22608:13
  assign _T_144 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22609:13
  mult mult_inst229 (	// matmul/matmul-hw.mlir:22610:28
    .a      (A_reg_bank229_p0_rd_data),	// matmul/matmul-hw.mlir:12444:33
    .b      (_T_2548),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst229_result)
  );
  assign _T_143 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22611:13
  assign a_i_k_5_i_j_14 = A_reg_bank229_p0_rd_data;	// matmul/matmul-hw.mlir:12444:33, :22613:5
  //PROBE: a_i_k_5_i_j_14	// matmul/matmul-hw.mlir:22614:5
  assign b_i_k_5_i_j_14 = _T_2548;	// matmul/matmul-hw.mlir:22616:5
  //PROBE: b_i_k_5_i_j_14	// matmul/matmul-hw.mlir:22617:5
  assign c_prev_i_k_5_i_j_14 = C_reg_bank5_p0_rd_data_2210;	// matmul/matmul-hw.mlir:22444:36, :22619:5
  //PROBE: c_prev_i_k_5_i_j_14	// matmul/matmul-hw.mlir:22620:5
  assign tk_i_k_5_i_j_14 = _T_2902;	// matmul/matmul-hw.mlir:22622:5
  //PROBE: tk_i_k_5_i_j_14	// matmul/matmul-hw.mlir:22623:5
  wire [31:0] _T_3948 = mult_inst229_result + C_reg_bank5_p0_rd_data_2210;	// matmul/matmul-hw.mlir:22444:36, :22610:28, :22624:13
  assign c_i_k_5_i_j_14 = _T_3948;	// matmul/matmul-hw.mlir:22626:5
  //PROBE: c_i_k_5_i_j_14	// matmul/matmul-hw.mlir:22627:5
  assign _T_142 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22628:13
  assign _T_141 = _T_2922 ? _T_3948 : 32'bx;	// matmul/matmul-hw.mlir:8176:18, :22629:13
  localparam [3:0] _T_3950 = 4'h0;	// matmul/matmul-hw.mlir:22632:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22633:5
    if (rst)	// matmul/matmul-hw.mlir:22633:5
      i_k_next_3949 <= _T_3950;	// matmul/matmul-hw.mlir:22636:7
    else	// matmul/matmul-hw.mlir:22633:5
      i_k_next_3949 <= i_k_next_3946;	// matmul/matmul-hw.mlir:22601:13, :22634:7
  end // always @(posedge)
  assign _T_140 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22638:13
  assign _T_139 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22639:13
  mult mult_inst230 (	// matmul/matmul-hw.mlir:22640:28
    .a      (A_reg_bank230_p0_rd_data),	// matmul/matmul-hw.mlir:12445:33
    .b      (_T_2564),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst230_result)
  );
  assign _T_138 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22641:13
  assign a_i_k_6_i_j_14 = A_reg_bank230_p0_rd_data;	// matmul/matmul-hw.mlir:12445:33, :22643:5
  //PROBE: a_i_k_6_i_j_14	// matmul/matmul-hw.mlir:22644:5
  assign b_i_k_6_i_j_14 = _T_2564;	// matmul/matmul-hw.mlir:22646:5
  //PROBE: b_i_k_6_i_j_14	// matmul/matmul-hw.mlir:22647:5
  assign c_prev_i_k_6_i_j_14 = C_reg_bank6_p0_rd_data_2209;	// matmul/matmul-hw.mlir:22445:36, :22649:5
  //PROBE: c_prev_i_k_6_i_j_14	// matmul/matmul-hw.mlir:22650:5
  assign tk_i_k_6_i_j_14 = _T_2907;	// matmul/matmul-hw.mlir:22652:5
  //PROBE: tk_i_k_6_i_j_14	// matmul/matmul-hw.mlir:22653:5
  wire [31:0] _T_3951 = mult_inst230_result + C_reg_bank6_p0_rd_data_2209;	// matmul/matmul-hw.mlir:22445:36, :22640:28, :22654:13
  assign c_i_k_6_i_j_14 = _T_3951;	// matmul/matmul-hw.mlir:22656:5
  //PROBE: c_i_k_6_i_j_14	// matmul/matmul-hw.mlir:22657:5
  assign _T_137 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22658:13
  assign _T_136 = _T_2927 ? _T_3951 : 32'bx;	// matmul/matmul-hw.mlir:8171:18, :22659:13
  localparam [3:0] _T_3953 = 4'h0;	// matmul/matmul-hw.mlir:22662:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22663:5
    if (rst)	// matmul/matmul-hw.mlir:22663:5
      i_k_next_3952 <= _T_3953;	// matmul/matmul-hw.mlir:22666:7
    else	// matmul/matmul-hw.mlir:22663:5
      i_k_next_3952 <= i_k_next_3949;	// matmul/matmul-hw.mlir:22631:13, :22664:7
  end // always @(posedge)
  assign _T_135 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22668:13
  assign _T_134 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22669:13
  mult mult_inst231 (	// matmul/matmul-hw.mlir:22670:28
    .a      (A_reg_bank231_p0_rd_data),	// matmul/matmul-hw.mlir:12446:33
    .b      (_T_2580),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst231_result)
  );
  assign _T_133 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22671:13
  assign a_i_k_7_i_j_14 = A_reg_bank231_p0_rd_data;	// matmul/matmul-hw.mlir:12446:33, :22673:5
  //PROBE: a_i_k_7_i_j_14	// matmul/matmul-hw.mlir:22674:5
  assign b_i_k_7_i_j_14 = _T_2580;	// matmul/matmul-hw.mlir:22676:5
  //PROBE: b_i_k_7_i_j_14	// matmul/matmul-hw.mlir:22677:5
  assign c_prev_i_k_7_i_j_14 = C_reg_bank7_p0_rd_data_2208;	// matmul/matmul-hw.mlir:22446:36, :22679:5
  //PROBE: c_prev_i_k_7_i_j_14	// matmul/matmul-hw.mlir:22680:5
  assign tk_i_k_7_i_j_14 = _T_2912;	// matmul/matmul-hw.mlir:22682:5
  //PROBE: tk_i_k_7_i_j_14	// matmul/matmul-hw.mlir:22683:5
  wire [31:0] _T_3954 = mult_inst231_result + C_reg_bank7_p0_rd_data_2208;	// matmul/matmul-hw.mlir:22446:36, :22670:28, :22684:13
  assign c_i_k_7_i_j_14 = _T_3954;	// matmul/matmul-hw.mlir:22686:5
  //PROBE: c_i_k_7_i_j_14	// matmul/matmul-hw.mlir:22687:5
  assign _T_132 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22688:13
  assign _T_131 = _T_2932 ? _T_3954 : 32'bx;	// matmul/matmul-hw.mlir:8166:18, :22689:13
  localparam [3:0] _T_3956 = 4'h0;	// matmul/matmul-hw.mlir:22692:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22693:5
    if (rst)	// matmul/matmul-hw.mlir:22693:5
      i_k_next_3955 <= _T_3956;	// matmul/matmul-hw.mlir:22696:7
    else	// matmul/matmul-hw.mlir:22693:5
      i_k_next_3955 <= i_k_next_3952;	// matmul/matmul-hw.mlir:22661:13, :22694:7
  end // always @(posedge)
  assign _T_130 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22698:13
  assign _T_129 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22699:13
  mult mult_inst232 (	// matmul/matmul-hw.mlir:22700:28
    .a      (A_reg_bank232_p0_rd_data),	// matmul/matmul-hw.mlir:12447:33
    .b      (_T_2596),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst232_result)
  );
  assign _T_128 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22701:13
  assign a_i_k_8_i_j_14 = A_reg_bank232_p0_rd_data;	// matmul/matmul-hw.mlir:12447:33, :22703:5
  //PROBE: a_i_k_8_i_j_14	// matmul/matmul-hw.mlir:22704:5
  assign b_i_k_8_i_j_14 = _T_2596;	// matmul/matmul-hw.mlir:22706:5
  //PROBE: b_i_k_8_i_j_14	// matmul/matmul-hw.mlir:22707:5
  assign c_prev_i_k_8_i_j_14 = C_reg_bank8_p0_rd_data_2207;	// matmul/matmul-hw.mlir:22447:36, :22709:5
  //PROBE: c_prev_i_k_8_i_j_14	// matmul/matmul-hw.mlir:22710:5
  assign tk_i_k_8_i_j_14 = _T_2917;	// matmul/matmul-hw.mlir:22712:5
  //PROBE: tk_i_k_8_i_j_14	// matmul/matmul-hw.mlir:22713:5
  wire [31:0] _T_3957 = mult_inst232_result + C_reg_bank8_p0_rd_data_2207;	// matmul/matmul-hw.mlir:22447:36, :22700:28, :22714:13
  assign c_i_k_8_i_j_14 = _T_3957;	// matmul/matmul-hw.mlir:22716:5
  //PROBE: c_i_k_8_i_j_14	// matmul/matmul-hw.mlir:22717:5
  assign _T_127 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22718:13
  assign _T_126 = _T_2937 ? _T_3957 : 32'bx;	// matmul/matmul-hw.mlir:8161:18, :22719:13
  localparam [3:0] _T_3959 = 4'h0;	// matmul/matmul-hw.mlir:22722:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22723:5
    if (rst)	// matmul/matmul-hw.mlir:22723:5
      i_k_next_3958 <= _T_3959;	// matmul/matmul-hw.mlir:22726:7
    else	// matmul/matmul-hw.mlir:22723:5
      i_k_next_3958 <= i_k_next_3955;	// matmul/matmul-hw.mlir:22691:13, :22724:7
  end // always @(posedge)
  assign _T_125 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22728:13
  assign _T_124 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22729:13
  mult mult_inst233 (	// matmul/matmul-hw.mlir:22730:28
    .a      (A_reg_bank233_p0_rd_data),	// matmul/matmul-hw.mlir:12448:33
    .b      (_T_2612),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst233_result)
  );
  assign _T_123 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22731:13
  assign a_i_k_9_i_j_14 = A_reg_bank233_p0_rd_data;	// matmul/matmul-hw.mlir:12448:33, :22733:5
  //PROBE: a_i_k_9_i_j_14	// matmul/matmul-hw.mlir:22734:5
  assign b_i_k_9_i_j_14 = _T_2612;	// matmul/matmul-hw.mlir:22736:5
  //PROBE: b_i_k_9_i_j_14	// matmul/matmul-hw.mlir:22737:5
  assign c_prev_i_k_9_i_j_14 = C_reg_bank9_p0_rd_data_2206;	// matmul/matmul-hw.mlir:22448:36, :22739:5
  //PROBE: c_prev_i_k_9_i_j_14	// matmul/matmul-hw.mlir:22740:5
  assign tk_i_k_9_i_j_14 = _T_2922;	// matmul/matmul-hw.mlir:22742:5
  //PROBE: tk_i_k_9_i_j_14	// matmul/matmul-hw.mlir:22743:5
  wire [31:0] _T_3960 = mult_inst233_result + C_reg_bank9_p0_rd_data_2206;	// matmul/matmul-hw.mlir:22448:36, :22730:28, :22744:13
  assign c_i_k_9_i_j_14 = _T_3960;	// matmul/matmul-hw.mlir:22746:5
  //PROBE: c_i_k_9_i_j_14	// matmul/matmul-hw.mlir:22747:5
  assign _T_122 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22748:13
  assign _T_121 = _T_2942 ? _T_3960 : 32'bx;	// matmul/matmul-hw.mlir:8156:18, :22749:13
  localparam [3:0] _T_3962 = 4'h0;	// matmul/matmul-hw.mlir:22752:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22753:5
    if (rst)	// matmul/matmul-hw.mlir:22753:5
      i_k_next_3961 <= _T_3962;	// matmul/matmul-hw.mlir:22756:7
    else	// matmul/matmul-hw.mlir:22753:5
      i_k_next_3961 <= i_k_next_3958;	// matmul/matmul-hw.mlir:22721:13, :22754:7
  end // always @(posedge)
  assign _T_120 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22758:13
  assign _T_119 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22759:13
  mult mult_inst234 (	// matmul/matmul-hw.mlir:22760:28
    .a      (A_reg_bank234_p0_rd_data),	// matmul/matmul-hw.mlir:12449:33
    .b      (_T_2628),
    .t      (_T_2937),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst234_result)
  );
  assign _T_118 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22761:13
  assign a_i_k_10_i_j_14 = A_reg_bank234_p0_rd_data;	// matmul/matmul-hw.mlir:12449:33, :22763:5
  //PROBE: a_i_k_10_i_j_14	// matmul/matmul-hw.mlir:22764:5
  assign b_i_k_10_i_j_14 = _T_2628;	// matmul/matmul-hw.mlir:22766:5
  //PROBE: b_i_k_10_i_j_14	// matmul/matmul-hw.mlir:22767:5
  assign c_prev_i_k_10_i_j_14 = C_reg_bank10_p0_rd_data_2205;	// matmul/matmul-hw.mlir:22449:37, :22769:5
  //PROBE: c_prev_i_k_10_i_j_14	// matmul/matmul-hw.mlir:22770:5
  assign tk_i_k_10_i_j_14 = _T_2927;	// matmul/matmul-hw.mlir:22772:5
  //PROBE: tk_i_k_10_i_j_14	// matmul/matmul-hw.mlir:22773:5
  wire [31:0] _T_3963 = mult_inst234_result + C_reg_bank10_p0_rd_data_2205;	// matmul/matmul-hw.mlir:22449:37, :22760:28, :22774:13
  assign c_i_k_10_i_j_14 = _T_3963;	// matmul/matmul-hw.mlir:22776:5
  //PROBE: c_i_k_10_i_j_14	// matmul/matmul-hw.mlir:22777:5
  assign _T_117 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22778:13
  assign _T_116 = _T_2947 ? _T_3963 : 32'bx;	// matmul/matmul-hw.mlir:8151:18, :22779:13
  localparam [3:0] _T_3965 = 4'h0;	// matmul/matmul-hw.mlir:22782:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22783:5
    if (rst)	// matmul/matmul-hw.mlir:22783:5
      i_k_next_3964 <= _T_3965;	// matmul/matmul-hw.mlir:22786:7
    else	// matmul/matmul-hw.mlir:22783:5
      i_k_next_3964 <= i_k_next_3961;	// matmul/matmul-hw.mlir:22751:13, :22784:7
  end // always @(posedge)
  assign _T_115 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22788:13
  assign _T_114 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22789:13
  mult mult_inst235 (	// matmul/matmul-hw.mlir:22790:28
    .a      (A_reg_bank235_p0_rd_data),	// matmul/matmul-hw.mlir:12450:33
    .b      (_T_2644),
    .t      (_T_2942),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst235_result)
  );
  assign _T_113 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22791:13
  assign a_i_k_11_i_j_14 = A_reg_bank235_p0_rd_data;	// matmul/matmul-hw.mlir:12450:33, :22793:5
  //PROBE: a_i_k_11_i_j_14	// matmul/matmul-hw.mlir:22794:5
  assign b_i_k_11_i_j_14 = _T_2644;	// matmul/matmul-hw.mlir:22796:5
  //PROBE: b_i_k_11_i_j_14	// matmul/matmul-hw.mlir:22797:5
  assign c_prev_i_k_11_i_j_14 = C_reg_bank11_p0_rd_data_2204;	// matmul/matmul-hw.mlir:22450:37, :22799:5
  //PROBE: c_prev_i_k_11_i_j_14	// matmul/matmul-hw.mlir:22800:5
  assign tk_i_k_11_i_j_14 = _T_2932;	// matmul/matmul-hw.mlir:22802:5
  //PROBE: tk_i_k_11_i_j_14	// matmul/matmul-hw.mlir:22803:5
  wire [31:0] _T_3966 = mult_inst235_result + C_reg_bank11_p0_rd_data_2204;	// matmul/matmul-hw.mlir:22450:37, :22790:28, :22804:13
  assign c_i_k_11_i_j_14 = _T_3966;	// matmul/matmul-hw.mlir:22806:5
  //PROBE: c_i_k_11_i_j_14	// matmul/matmul-hw.mlir:22807:5
  assign _T_112 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22808:13
  assign _T_111 = _T_2952 ? _T_3966 : 32'bx;	// matmul/matmul-hw.mlir:8146:18, :22809:13
  localparam [3:0] _T_3968 = 4'h0;	// matmul/matmul-hw.mlir:22812:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22813:5
    if (rst)	// matmul/matmul-hw.mlir:22813:5
      i_k_next_3967 <= _T_3968;	// matmul/matmul-hw.mlir:22816:7
    else	// matmul/matmul-hw.mlir:22813:5
      i_k_next_3967 <= i_k_next_3964;	// matmul/matmul-hw.mlir:22781:13, :22814:7
  end // always @(posedge)
  assign _T_110 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22818:13
  assign _T_109 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22819:13
  mult mult_inst236 (	// matmul/matmul-hw.mlir:22820:28
    .a      (A_reg_bank236_p0_rd_data),	// matmul/matmul-hw.mlir:12451:33
    .b      (_T_2660),
    .t      (_T_2947),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst236_result)
  );
  assign _T_108 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22821:13
  assign a_i_k_12_i_j_14 = A_reg_bank236_p0_rd_data;	// matmul/matmul-hw.mlir:12451:33, :22823:5
  //PROBE: a_i_k_12_i_j_14	// matmul/matmul-hw.mlir:22824:5
  assign b_i_k_12_i_j_14 = _T_2660;	// matmul/matmul-hw.mlir:22826:5
  //PROBE: b_i_k_12_i_j_14	// matmul/matmul-hw.mlir:22827:5
  assign c_prev_i_k_12_i_j_14 = C_reg_bank12_p0_rd_data_2203;	// matmul/matmul-hw.mlir:22451:37, :22829:5
  //PROBE: c_prev_i_k_12_i_j_14	// matmul/matmul-hw.mlir:22830:5
  assign tk_i_k_12_i_j_14 = _T_2937;	// matmul/matmul-hw.mlir:22832:5
  //PROBE: tk_i_k_12_i_j_14	// matmul/matmul-hw.mlir:22833:5
  wire [31:0] _T_3969 = mult_inst236_result + C_reg_bank12_p0_rd_data_2203;	// matmul/matmul-hw.mlir:22451:37, :22820:28, :22834:13
  assign c_i_k_12_i_j_14 = _T_3969;	// matmul/matmul-hw.mlir:22836:5
  //PROBE: c_i_k_12_i_j_14	// matmul/matmul-hw.mlir:22837:5
  assign _T_107 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22838:13
  assign _T_106 = _T_2957 ? _T_3969 : 32'bx;	// matmul/matmul-hw.mlir:8141:18, :22839:13
  localparam [3:0] _T_3971 = 4'h0;	// matmul/matmul-hw.mlir:22842:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22843:5
    if (rst)	// matmul/matmul-hw.mlir:22843:5
      i_k_next_3970 <= _T_3971;	// matmul/matmul-hw.mlir:22846:7
    else	// matmul/matmul-hw.mlir:22843:5
      i_k_next_3970 <= i_k_next_3967;	// matmul/matmul-hw.mlir:22811:13, :22844:7
  end // always @(posedge)
  assign _T_105 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22848:13
  assign _T_104 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22849:13
  mult mult_inst237 (	// matmul/matmul-hw.mlir:22850:28
    .a      (A_reg_bank237_p0_rd_data),	// matmul/matmul-hw.mlir:12452:33
    .b      (_T_2676),
    .t      (_T_2952),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst237_result)
  );
  assign _T_103 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22851:13
  assign a_i_k_13_i_j_14 = A_reg_bank237_p0_rd_data;	// matmul/matmul-hw.mlir:12452:33, :22853:5
  //PROBE: a_i_k_13_i_j_14	// matmul/matmul-hw.mlir:22854:5
  assign b_i_k_13_i_j_14 = _T_2676;	// matmul/matmul-hw.mlir:22856:5
  //PROBE: b_i_k_13_i_j_14	// matmul/matmul-hw.mlir:22857:5
  assign c_prev_i_k_13_i_j_14 = C_reg_bank13_p0_rd_data_2202;	// matmul/matmul-hw.mlir:22452:37, :22859:5
  //PROBE: c_prev_i_k_13_i_j_14	// matmul/matmul-hw.mlir:22860:5
  assign tk_i_k_13_i_j_14 = _T_2942;	// matmul/matmul-hw.mlir:22862:5
  //PROBE: tk_i_k_13_i_j_14	// matmul/matmul-hw.mlir:22863:5
  wire [31:0] _T_3972 = mult_inst237_result + C_reg_bank13_p0_rd_data_2202;	// matmul/matmul-hw.mlir:22452:37, :22850:28, :22864:13
  assign c_i_k_13_i_j_14 = _T_3972;	// matmul/matmul-hw.mlir:22866:5
  //PROBE: c_i_k_13_i_j_14	// matmul/matmul-hw.mlir:22867:5
  assign _T_102 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22868:13
  assign _T_101 = _T_2962 ? _T_3972 : 32'bx;	// matmul/matmul-hw.mlir:8136:18, :22869:13
  localparam [3:0] _T_3974 = 4'h0;	// matmul/matmul-hw.mlir:22872:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22873:5
    if (rst)	// matmul/matmul-hw.mlir:22873:5
      i_k_next_3973 <= _T_3974;	// matmul/matmul-hw.mlir:22876:7
    else	// matmul/matmul-hw.mlir:22873:5
      i_k_next_3973 <= i_k_next_3970;	// matmul/matmul-hw.mlir:22841:13, :22874:7
  end // always @(posedge)
  assign _T_100 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22878:13
  assign _T_99 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22879:13
  mult mult_inst238 (	// matmul/matmul-hw.mlir:22880:28
    .a      (A_reg_bank238_p0_rd_data),	// matmul/matmul-hw.mlir:12453:33
    .b      (_T_2692),
    .t      (_T_2957),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst238_result)
  );
  assign _T_98 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22881:13
  assign a_i_k_14_i_j_14 = A_reg_bank238_p0_rd_data;	// matmul/matmul-hw.mlir:12453:33, :22883:5
  //PROBE: a_i_k_14_i_j_14	// matmul/matmul-hw.mlir:22884:5
  assign b_i_k_14_i_j_14 = _T_2692;	// matmul/matmul-hw.mlir:22886:5
  //PROBE: b_i_k_14_i_j_14	// matmul/matmul-hw.mlir:22887:5
  assign c_prev_i_k_14_i_j_14 = C_reg_bank14_p0_rd_data_2201;	// matmul/matmul-hw.mlir:22453:37, :22889:5
  //PROBE: c_prev_i_k_14_i_j_14	// matmul/matmul-hw.mlir:22890:5
  assign tk_i_k_14_i_j_14 = _T_2947;	// matmul/matmul-hw.mlir:22892:5
  //PROBE: tk_i_k_14_i_j_14	// matmul/matmul-hw.mlir:22893:5
  wire [31:0] _T_3975 = mult_inst238_result + C_reg_bank14_p0_rd_data_2201;	// matmul/matmul-hw.mlir:22453:37, :22880:28, :22894:13
  assign c_i_k_14_i_j_14 = _T_3975;	// matmul/matmul-hw.mlir:22896:5
  //PROBE: c_i_k_14_i_j_14	// matmul/matmul-hw.mlir:22897:5
  assign _T_97 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22898:13
  assign _T_96 = _T_3833 ? _T_3975 : 32'bx;	// matmul/matmul-hw.mlir:8131:18, :22899:13
  localparam [3:0] _T_3977 = 4'h0;	// matmul/matmul-hw.mlir:22902:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22903:5
    if (rst)	// matmul/matmul-hw.mlir:22903:5
      i_k_next_3976 <= _T_3977;	// matmul/matmul-hw.mlir:22906:7
    else	// matmul/matmul-hw.mlir:22903:5
      i_k_next_3976 <= i_k_next_3973;	// matmul/matmul-hw.mlir:22871:13, :22904:7
  end // always @(posedge)
  assign _T_95 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22908:13
  assign _T_94 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22909:13
  mult mult_inst239 (	// matmul/matmul-hw.mlir:22910:28
    .a      (A_reg_bank239_p0_rd_data),	// matmul/matmul-hw.mlir:12454:33
    .b      (_T_2708),
    .t      (_T_2962),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst239_result)
  );
  assign _T_93 = _T_3909 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22911:13
  assign a_i_k_15_i_j_14 = A_reg_bank239_p0_rd_data;	// matmul/matmul-hw.mlir:12454:33, :22913:5
  //PROBE: a_i_k_15_i_j_14	// matmul/matmul-hw.mlir:22914:5
  assign b_i_k_15_i_j_14 = _T_2708;	// matmul/matmul-hw.mlir:22916:5
  //PROBE: b_i_k_15_i_j_14	// matmul/matmul-hw.mlir:22917:5
  assign c_prev_i_k_15_i_j_14 = C_reg_bank15_p0_rd_data_2200;	// matmul/matmul-hw.mlir:22454:37, :22919:5
  //PROBE: c_prev_i_k_15_i_j_14	// matmul/matmul-hw.mlir:22920:5
  assign tk_i_k_15_i_j_14 = _T_2952;	// matmul/matmul-hw.mlir:22922:5
  //PROBE: tk_i_k_15_i_j_14	// matmul/matmul-hw.mlir:22923:5
  wire [31:0] _T_3978 = mult_inst239_result + C_reg_bank15_p0_rd_data_2200;	// matmul/matmul-hw.mlir:22454:37, :22910:28, :22924:13
  assign c_i_k_15_i_j_14 = _T_3978;	// matmul/matmul-hw.mlir:22926:5
  //PROBE: c_i_k_15_i_j_14	// matmul/matmul-hw.mlir:22927:5
  assign _T_92 = _T_3909 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22928:13
  assign _T_91 = _T_3909 ? _T_3978 : 32'bx;	// matmul/matmul-hw.mlir:8126:18, :22929:13
  localparam [3:0] _T_3980 = 4'h0;	// matmul/matmul-hw.mlir:22932:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22933:5
    if (rst)	// matmul/matmul-hw.mlir:22933:5
      i_k_next_3979 <= _T_3980;	// matmul/matmul-hw.mlir:22936:7
    else	// matmul/matmul-hw.mlir:22933:5
      i_k_next_3979 <= i_k_next_3976;	// matmul/matmul-hw.mlir:22901:13, :22934:7
  end // always @(posedge)
  wire [33:0] _T_3982 = _T_3981;	// matmul/matmul-hw.mlir:22939:13
  wire [33:0] _T_3983 = {_T_3982[6'h0+:33], {{_T_2712}}};	// matmul/matmul-hw.mlir:22940:19, :22941:13, :22942:13, :22943:13
  wire [33:0] _T_3984 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:22944:19, :22945:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22946:5
    if (rst)	// matmul/matmul-hw.mlir:22946:5
      _T_3981 <= _T_3984;	// matmul/matmul-hw.mlir:22949:7
    else	// matmul/matmul-hw.mlir:22946:5
      _T_3981 <= _T_3983;	// matmul/matmul-hw.mlir:22947:7
  end // always @(posedge)
  wire _T_3985 = _T_3981[6'h21];	// matmul/matmul-hw.mlir:22939:13, :22951:16, :22952:13
  assign _T_90 = _T_3985 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22953:13
  wire [3:0][3:0] _T_3987 = i_delayed_3986;	// matmul/matmul-hw.mlir:22955:13
  wire [3:0][3:0] _T_3988 = {_T_3987[2'h0+:3], {{i_k_next_3979}}};	// matmul/matmul-hw.mlir:22931:13, :22956:19, :22957:13, :22958:13, :22959:13
  wire [3:0][3:0] _T_3989 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:22960:19, :22961:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22962:5
    if (rst)	// matmul/matmul-hw.mlir:22962:5
      i_delayed_3986 <= _T_3989;	// matmul/matmul-hw.mlir:22965:7
    else	// matmul/matmul-hw.mlir:22962:5
      i_delayed_3986 <= _T_3988;	// matmul/matmul-hw.mlir:22963:7
  end // always @(posedge)
  assign _T_89 = _T_3985 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22969:13
  assign _T_88 = _T_3985 ? i_delayed_3986[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8123:17, :22955:13, :22967:20, :22968:13, :22970:13
  assign _T_87 = _T_3985 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :22971:13
  assign _T_86 = _T_3985 ? C_reg_bank16_p0_rd_data_2199 : 32'bx;	// matmul/matmul-hw.mlir:8121:18, :22455:37, :22972:13
  localparam [3:0] _T_3991 = 4'h0;	// matmul/matmul-hw.mlir:22975:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:22976:5
    if (rst)	// matmul/matmul-hw.mlir:22976:5
      i_j_next_3990 <= _T_3991;	// matmul/matmul-hw.mlir:22979:7
    else	// matmul/matmul-hw.mlir:22976:5
      i_j_next_3990 <= i_j_next_3914;	// matmul/matmul-hw.mlir:22364:13, :22977:7
  end // always @(posedge)
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank0_3992 (	// matmul/matmul-hw.mlir:23049:36
    .p0_rd_en   (_T_81),	// matmul/matmul-hw.mlir:23071:13
    .p1_wr_en   (_T_85),	// matmul/matmul-hw.mlir:23066:13
    .p1_wr_data (_T_84),	// matmul/matmul-hw.mlir:23067:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank0_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank1_3993 (	// matmul/matmul-hw.mlir:23050:36
    .p0_rd_en   (_T_76),	// matmul/matmul-hw.mlir:23101:13
    .p1_wr_en   (_T_80),	// matmul/matmul-hw.mlir:23088:13
    .p1_wr_data (_T_79),	// matmul/matmul-hw.mlir:23089:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank1_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank2_3994 (	// matmul/matmul-hw.mlir:23051:36
    .p0_rd_en   (_T_71),	// matmul/matmul-hw.mlir:23131:13
    .p1_wr_en   (_T_75),	// matmul/matmul-hw.mlir:23118:13
    .p1_wr_data (_T_74),	// matmul/matmul-hw.mlir:23119:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank2_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank3_3995 (	// matmul/matmul-hw.mlir:23052:36
    .p0_rd_en   (_T_66),	// matmul/matmul-hw.mlir:23161:13
    .p1_wr_en   (_T_70),	// matmul/matmul-hw.mlir:23148:13
    .p1_wr_data (_T_69),	// matmul/matmul-hw.mlir:23149:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank3_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank4_3996 (	// matmul/matmul-hw.mlir:23053:36
    .p0_rd_en   (_T_61),	// matmul/matmul-hw.mlir:23191:13
    .p1_wr_en   (_T_65),	// matmul/matmul-hw.mlir:23178:13
    .p1_wr_data (_T_64),	// matmul/matmul-hw.mlir:23179:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank4_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank5_3997 (	// matmul/matmul-hw.mlir:23054:36
    .p0_rd_en   (_T_56),	// matmul/matmul-hw.mlir:23221:13
    .p1_wr_en   (_T_60),	// matmul/matmul-hw.mlir:23208:13
    .p1_wr_data (_T_59),	// matmul/matmul-hw.mlir:23209:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank5_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank6_3998 (	// matmul/matmul-hw.mlir:23055:36
    .p0_rd_en   (_T_51),	// matmul/matmul-hw.mlir:23251:13
    .p1_wr_en   (_T_55),	// matmul/matmul-hw.mlir:23238:13
    .p1_wr_data (_T_54),	// matmul/matmul-hw.mlir:23239:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank6_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank7_3999 (	// matmul/matmul-hw.mlir:23056:36
    .p0_rd_en   (_T_46),	// matmul/matmul-hw.mlir:23281:13
    .p1_wr_en   (_T_50),	// matmul/matmul-hw.mlir:23268:13
    .p1_wr_data (_T_49),	// matmul/matmul-hw.mlir:23269:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank7_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank8_4000 (	// matmul/matmul-hw.mlir:23057:36
    .p0_rd_en   (_T_41),	// matmul/matmul-hw.mlir:23311:13
    .p1_wr_en   (_T_45),	// matmul/matmul-hw.mlir:23298:13
    .p1_wr_data (_T_44),	// matmul/matmul-hw.mlir:23299:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank8_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank9_4001 (	// matmul/matmul-hw.mlir:23058:36
    .p0_rd_en   (_T_36),	// matmul/matmul-hw.mlir:23341:13
    .p1_wr_en   (_T_40),	// matmul/matmul-hw.mlir:23328:13
    .p1_wr_data (_T_39),	// matmul/matmul-hw.mlir:23329:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank9_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank10_4002 (	// matmul/matmul-hw.mlir:23059:37
    .p0_rd_en   (_T_31),	// matmul/matmul-hw.mlir:23371:13
    .p1_wr_en   (_T_35),	// matmul/matmul-hw.mlir:23358:13
    .p1_wr_data (_T_34),	// matmul/matmul-hw.mlir:23359:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank10_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank11_4003 (	// matmul/matmul-hw.mlir:23060:37
    .p0_rd_en   (_T_26),	// matmul/matmul-hw.mlir:23401:13
    .p1_wr_en   (_T_30),	// matmul/matmul-hw.mlir:23388:13
    .p1_wr_data (_T_29),	// matmul/matmul-hw.mlir:23389:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank11_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank12_4004 (	// matmul/matmul-hw.mlir:23061:37
    .p0_rd_en   (_T_21),	// matmul/matmul-hw.mlir:23431:13
    .p1_wr_en   (_T_25),	// matmul/matmul-hw.mlir:23418:13
    .p1_wr_data (_T_24),	// matmul/matmul-hw.mlir:23419:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank12_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank13_4005 (	// matmul/matmul-hw.mlir:23062:37
    .p0_rd_en   (_T_16),	// matmul/matmul-hw.mlir:23461:13
    .p1_wr_en   (_T_20),	// matmul/matmul-hw.mlir:23448:13
    .p1_wr_data (_T_19),	// matmul/matmul-hw.mlir:23449:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank13_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank14_4006 (	// matmul/matmul-hw.mlir:23063:37
    .p0_rd_en   (_T_11),	// matmul/matmul-hw.mlir:23491:13
    .p1_wr_en   (_T_15),	// matmul/matmul-hw.mlir:23478:13
    .p1_wr_data (_T_14),	// matmul/matmul-hw.mlir:23479:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank14_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank15_4007 (	// matmul/matmul-hw.mlir:23064:37
    .p0_rd_en   (_T_6),	// matmul/matmul-hw.mlir:23521:13
    .p1_wr_en   (_T_10),	// matmul/matmul-hw.mlir:23508:13
    .p1_wr_data (_T_9),	// matmul/matmul-hw.mlir:23509:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank15_p0_rd_data)
  );
  reg_r0_w1 #(
    .ELEMENT_WIDTH(64'd32)
  ) C_reg_bank16_4008 (	// matmul/matmul-hw.mlir:23065:37
    .p0_rd_en   (_T_3),	// matmul/matmul-hw.mlir:23563:13
    .p1_wr_en   (_T_5),	// matmul/matmul-hw.mlir:23538:13
    .p1_wr_data (_T_4),	// matmul/matmul-hw.mlir:23539:13
    .t          (_T_2712),
    .clk        (clk),
    .rst        (rst),
    .p0_rd_data (C_reg_bank16_p0_rd_data)
  );
  assign _T_85 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23066:13
  assign _T_84 = _T_2897 ? 32'h0 : 32'bx;	// matmul/matmul-hw.mlir:8028:15, :8119:18, :23067:13
  assign _T_83 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23068:13
  assign _T_82 = _T_2892 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23069:13
  mult mult_inst240 (	// matmul/matmul-hw.mlir:23070:28
    .a      (A_reg_bank240_p0_rd_data),	// matmul/matmul-hw.mlir:12455:33
    .b      (_T_2469),
    .t      (_T_2892),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst240_result)
  );
  assign _T_81 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23071:13
  assign a_i_k_0_i_j_15 = A_reg_bank240_p0_rd_data;	// matmul/matmul-hw.mlir:12455:33, :23073:5
  //PROBE: a_i_k_0_i_j_15	// matmul/matmul-hw.mlir:23074:5
  assign b_i_k_0_i_j_15 = _T_2469;	// matmul/matmul-hw.mlir:23076:5
  //PROBE: b_i_k_0_i_j_15	// matmul/matmul-hw.mlir:23077:5
  assign c_prev_i_k_0_i_j_15 = C_reg_bank0_p0_rd_data;	// matmul/matmul-hw.mlir:23049:36, :23079:5
  //PROBE: c_prev_i_k_0_i_j_15	// matmul/matmul-hw.mlir:23080:5
  assign tk_i_k_0_i_j_15 = _T_2874;	// matmul/matmul-hw.mlir:23082:5
  //PROBE: tk_i_k_0_i_j_15	// matmul/matmul-hw.mlir:23083:5
  wire [31:0] _T_4009 = mult_inst240_result + C_reg_bank0_p0_rd_data;	// matmul/matmul-hw.mlir:23049:36, :23070:28, :23084:13
  assign c_i_k_0_i_j_15 = _T_4009;	// matmul/matmul-hw.mlir:23086:5
  //PROBE: c_i_k_0_i_j_15	// matmul/matmul-hw.mlir:23087:5
  assign _T_80 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23088:13
  assign _T_79 = _T_2902 ? _T_4009 : 32'bx;	// matmul/matmul-hw.mlir:8114:18, :23089:13
  localparam [3:0] _T_4011 = 4'h0;	// matmul/matmul-hw.mlir:23092:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23093:5
    if (rst)	// matmul/matmul-hw.mlir:23093:5
      i_k_next_4010 <= _T_4011;	// matmul/matmul-hw.mlir:23096:7
    else	// matmul/matmul-hw.mlir:23093:5
      i_k_next_4010 <= i_j_next_3990;	// matmul/matmul-hw.mlir:22974:13, :23094:7
  end // always @(posedge)
  assign _T_78 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23098:13
  assign _T_77 = _T_2897 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23099:13
  mult mult_inst241 (	// matmul/matmul-hw.mlir:23100:28
    .a      (A_reg_bank241_p0_rd_data),	// matmul/matmul-hw.mlir:12456:33
    .b      (_T_2485),
    .t      (_T_2897),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst241_result)
  );
  assign _T_76 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23101:13
  assign a_i_k_1_i_j_15 = A_reg_bank241_p0_rd_data;	// matmul/matmul-hw.mlir:12456:33, :23103:5
  //PROBE: a_i_k_1_i_j_15	// matmul/matmul-hw.mlir:23104:5
  assign b_i_k_1_i_j_15 = _T_2485;	// matmul/matmul-hw.mlir:23106:5
  //PROBE: b_i_k_1_i_j_15	// matmul/matmul-hw.mlir:23107:5
  assign c_prev_i_k_1_i_j_15 = C_reg_bank1_p0_rd_data;	// matmul/matmul-hw.mlir:23050:36, :23109:5
  //PROBE: c_prev_i_k_1_i_j_15	// matmul/matmul-hw.mlir:23110:5
  assign tk_i_k_1_i_j_15 = _T_2885;	// matmul/matmul-hw.mlir:23112:5
  //PROBE: tk_i_k_1_i_j_15	// matmul/matmul-hw.mlir:23113:5
  wire [31:0] _T_4012 = mult_inst241_result + C_reg_bank1_p0_rd_data;	// matmul/matmul-hw.mlir:23050:36, :23100:28, :23114:13
  assign c_i_k_1_i_j_15 = _T_4012;	// matmul/matmul-hw.mlir:23116:5
  //PROBE: c_i_k_1_i_j_15	// matmul/matmul-hw.mlir:23117:5
  assign _T_75 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23118:13
  assign _T_74 = _T_2907 ? _T_4012 : 32'bx;	// matmul/matmul-hw.mlir:8109:18, :23119:13
  localparam [3:0] _T_4014 = 4'h0;	// matmul/matmul-hw.mlir:23122:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23123:5
    if (rst)	// matmul/matmul-hw.mlir:23123:5
      i_k_next_4013 <= _T_4014;	// matmul/matmul-hw.mlir:23126:7
    else	// matmul/matmul-hw.mlir:23123:5
      i_k_next_4013 <= i_k_next_4010;	// matmul/matmul-hw.mlir:23091:13, :23124:7
  end // always @(posedge)
  assign _T_73 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23128:13
  assign _T_72 = _T_2902 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23129:13
  mult mult_inst242 (	// matmul/matmul-hw.mlir:23130:28
    .a      (A_reg_bank242_p0_rd_data),	// matmul/matmul-hw.mlir:12457:33
    .b      (_T_2501),
    .t      (_T_2902),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst242_result)
  );
  assign _T_71 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23131:13
  assign a_i_k_2_i_j_15 = A_reg_bank242_p0_rd_data;	// matmul/matmul-hw.mlir:12457:33, :23133:5
  //PROBE: a_i_k_2_i_j_15	// matmul/matmul-hw.mlir:23134:5
  assign b_i_k_2_i_j_15 = _T_2501;	// matmul/matmul-hw.mlir:23136:5
  //PROBE: b_i_k_2_i_j_15	// matmul/matmul-hw.mlir:23137:5
  assign c_prev_i_k_2_i_j_15 = C_reg_bank2_p0_rd_data;	// matmul/matmul-hw.mlir:23051:36, :23139:5
  //PROBE: c_prev_i_k_2_i_j_15	// matmul/matmul-hw.mlir:23140:5
  assign tk_i_k_2_i_j_15 = _T_2892;	// matmul/matmul-hw.mlir:23142:5
  //PROBE: tk_i_k_2_i_j_15	// matmul/matmul-hw.mlir:23143:5
  wire [31:0] _T_4015 = mult_inst242_result + C_reg_bank2_p0_rd_data;	// matmul/matmul-hw.mlir:23051:36, :23130:28, :23144:13
  assign c_i_k_2_i_j_15 = _T_4015;	// matmul/matmul-hw.mlir:23146:5
  //PROBE: c_i_k_2_i_j_15	// matmul/matmul-hw.mlir:23147:5
  assign _T_70 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23148:13
  assign _T_69 = _T_2912 ? _T_4015 : 32'bx;	// matmul/matmul-hw.mlir:8104:18, :23149:13
  localparam [3:0] _T_4017 = 4'h0;	// matmul/matmul-hw.mlir:23152:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23153:5
    if (rst)	// matmul/matmul-hw.mlir:23153:5
      i_k_next_4016 <= _T_4017;	// matmul/matmul-hw.mlir:23156:7
    else	// matmul/matmul-hw.mlir:23153:5
      i_k_next_4016 <= i_k_next_4013;	// matmul/matmul-hw.mlir:23121:13, :23154:7
  end // always @(posedge)
  assign _T_68 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23158:13
  assign _T_67 = _T_2907 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23159:13
  mult mult_inst243 (	// matmul/matmul-hw.mlir:23160:28
    .a      (A_reg_bank243_p0_rd_data),	// matmul/matmul-hw.mlir:12458:33
    .b      (_T_2517),
    .t      (_T_2907),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst243_result)
  );
  assign _T_66 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23161:13
  assign a_i_k_3_i_j_15 = A_reg_bank243_p0_rd_data;	// matmul/matmul-hw.mlir:12458:33, :23163:5
  //PROBE: a_i_k_3_i_j_15	// matmul/matmul-hw.mlir:23164:5
  assign b_i_k_3_i_j_15 = _T_2517;	// matmul/matmul-hw.mlir:23166:5
  //PROBE: b_i_k_3_i_j_15	// matmul/matmul-hw.mlir:23167:5
  assign c_prev_i_k_3_i_j_15 = C_reg_bank3_p0_rd_data;	// matmul/matmul-hw.mlir:23052:36, :23169:5
  //PROBE: c_prev_i_k_3_i_j_15	// matmul/matmul-hw.mlir:23170:5
  assign tk_i_k_3_i_j_15 = _T_2897;	// matmul/matmul-hw.mlir:23172:5
  //PROBE: tk_i_k_3_i_j_15	// matmul/matmul-hw.mlir:23173:5
  wire [31:0] _T_4018 = mult_inst243_result + C_reg_bank3_p0_rd_data;	// matmul/matmul-hw.mlir:23052:36, :23160:28, :23174:13
  assign c_i_k_3_i_j_15 = _T_4018;	// matmul/matmul-hw.mlir:23176:5
  //PROBE: c_i_k_3_i_j_15	// matmul/matmul-hw.mlir:23177:5
  assign _T_65 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23178:13
  assign _T_64 = _T_2917 ? _T_4018 : 32'bx;	// matmul/matmul-hw.mlir:8099:18, :23179:13
  localparam [3:0] _T_4020 = 4'h0;	// matmul/matmul-hw.mlir:23182:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23183:5
    if (rst)	// matmul/matmul-hw.mlir:23183:5
      i_k_next_4019 <= _T_4020;	// matmul/matmul-hw.mlir:23186:7
    else	// matmul/matmul-hw.mlir:23183:5
      i_k_next_4019 <= i_k_next_4016;	// matmul/matmul-hw.mlir:23151:13, :23184:7
  end // always @(posedge)
  assign _T_63 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23188:13
  assign _T_62 = _T_2912 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23189:13
  mult mult_inst244 (	// matmul/matmul-hw.mlir:23190:28
    .a      (A_reg_bank244_p0_rd_data),	// matmul/matmul-hw.mlir:12459:33
    .b      (_T_2533),
    .t      (_T_2912),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst244_result)
  );
  assign _T_61 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23191:13
  assign a_i_k_4_i_j_15 = A_reg_bank244_p0_rd_data;	// matmul/matmul-hw.mlir:12459:33, :23193:5
  //PROBE: a_i_k_4_i_j_15	// matmul/matmul-hw.mlir:23194:5
  assign b_i_k_4_i_j_15 = _T_2533;	// matmul/matmul-hw.mlir:23196:5
  //PROBE: b_i_k_4_i_j_15	// matmul/matmul-hw.mlir:23197:5
  assign c_prev_i_k_4_i_j_15 = C_reg_bank4_p0_rd_data;	// matmul/matmul-hw.mlir:23053:36, :23199:5
  //PROBE: c_prev_i_k_4_i_j_15	// matmul/matmul-hw.mlir:23200:5
  assign tk_i_k_4_i_j_15 = _T_2902;	// matmul/matmul-hw.mlir:23202:5
  //PROBE: tk_i_k_4_i_j_15	// matmul/matmul-hw.mlir:23203:5
  wire [31:0] _T_4021 = mult_inst244_result + C_reg_bank4_p0_rd_data;	// matmul/matmul-hw.mlir:23053:36, :23190:28, :23204:13
  assign c_i_k_4_i_j_15 = _T_4021;	// matmul/matmul-hw.mlir:23206:5
  //PROBE: c_i_k_4_i_j_15	// matmul/matmul-hw.mlir:23207:5
  assign _T_60 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23208:13
  assign _T_59 = _T_2922 ? _T_4021 : 32'bx;	// matmul/matmul-hw.mlir:8094:18, :23209:13
  localparam [3:0] _T_4023 = 4'h0;	// matmul/matmul-hw.mlir:23212:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23213:5
    if (rst)	// matmul/matmul-hw.mlir:23213:5
      i_k_next_4022 <= _T_4023;	// matmul/matmul-hw.mlir:23216:7
    else	// matmul/matmul-hw.mlir:23213:5
      i_k_next_4022 <= i_k_next_4019;	// matmul/matmul-hw.mlir:23181:13, :23214:7
  end // always @(posedge)
  assign _T_58 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23218:13
  assign _T_57 = _T_2917 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23219:13
  mult mult_inst245 (	// matmul/matmul-hw.mlir:23220:28
    .a      (A_reg_bank245_p0_rd_data),	// matmul/matmul-hw.mlir:12460:33
    .b      (_T_2549),
    .t      (_T_2917),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst245_result)
  );
  assign _T_56 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23221:13
  assign a_i_k_5_i_j_15 = A_reg_bank245_p0_rd_data;	// matmul/matmul-hw.mlir:12460:33, :23223:5
  //PROBE: a_i_k_5_i_j_15	// matmul/matmul-hw.mlir:23224:5
  assign b_i_k_5_i_j_15 = _T_2549;	// matmul/matmul-hw.mlir:23226:5
  //PROBE: b_i_k_5_i_j_15	// matmul/matmul-hw.mlir:23227:5
  assign c_prev_i_k_5_i_j_15 = C_reg_bank5_p0_rd_data;	// matmul/matmul-hw.mlir:23054:36, :23229:5
  //PROBE: c_prev_i_k_5_i_j_15	// matmul/matmul-hw.mlir:23230:5
  assign tk_i_k_5_i_j_15 = _T_2907;	// matmul/matmul-hw.mlir:23232:5
  //PROBE: tk_i_k_5_i_j_15	// matmul/matmul-hw.mlir:23233:5
  wire [31:0] _T_4024 = mult_inst245_result + C_reg_bank5_p0_rd_data;	// matmul/matmul-hw.mlir:23054:36, :23220:28, :23234:13
  assign c_i_k_5_i_j_15 = _T_4024;	// matmul/matmul-hw.mlir:23236:5
  //PROBE: c_i_k_5_i_j_15	// matmul/matmul-hw.mlir:23237:5
  assign _T_55 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23238:13
  assign _T_54 = _T_2927 ? _T_4024 : 32'bx;	// matmul/matmul-hw.mlir:8089:18, :23239:13
  localparam [3:0] _T_4026 = 4'h0;	// matmul/matmul-hw.mlir:23242:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23243:5
    if (rst)	// matmul/matmul-hw.mlir:23243:5
      i_k_next_4025 <= _T_4026;	// matmul/matmul-hw.mlir:23246:7
    else	// matmul/matmul-hw.mlir:23243:5
      i_k_next_4025 <= i_k_next_4022;	// matmul/matmul-hw.mlir:23211:13, :23244:7
  end // always @(posedge)
  assign _T_53 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23248:13
  assign _T_52 = _T_2922 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23249:13
  mult mult_inst246 (	// matmul/matmul-hw.mlir:23250:28
    .a      (A_reg_bank246_p0_rd_data),	// matmul/matmul-hw.mlir:12461:33
    .b      (_T_2565),
    .t      (_T_2922),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst246_result)
  );
  assign _T_51 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23251:13
  assign a_i_k_6_i_j_15 = A_reg_bank246_p0_rd_data;	// matmul/matmul-hw.mlir:12461:33, :23253:5
  //PROBE: a_i_k_6_i_j_15	// matmul/matmul-hw.mlir:23254:5
  assign b_i_k_6_i_j_15 = _T_2565;	// matmul/matmul-hw.mlir:23256:5
  //PROBE: b_i_k_6_i_j_15	// matmul/matmul-hw.mlir:23257:5
  assign c_prev_i_k_6_i_j_15 = C_reg_bank6_p0_rd_data;	// matmul/matmul-hw.mlir:23055:36, :23259:5
  //PROBE: c_prev_i_k_6_i_j_15	// matmul/matmul-hw.mlir:23260:5
  assign tk_i_k_6_i_j_15 = _T_2912;	// matmul/matmul-hw.mlir:23262:5
  //PROBE: tk_i_k_6_i_j_15	// matmul/matmul-hw.mlir:23263:5
  wire [31:0] _T_4027 = mult_inst246_result + C_reg_bank6_p0_rd_data;	// matmul/matmul-hw.mlir:23055:36, :23250:28, :23264:13
  assign c_i_k_6_i_j_15 = _T_4027;	// matmul/matmul-hw.mlir:23266:5
  //PROBE: c_i_k_6_i_j_15	// matmul/matmul-hw.mlir:23267:5
  assign _T_50 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23268:13
  assign _T_49 = _T_2932 ? _T_4027 : 32'bx;	// matmul/matmul-hw.mlir:8084:18, :23269:13
  localparam [3:0] _T_4029 = 4'h0;	// matmul/matmul-hw.mlir:23272:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23273:5
    if (rst)	// matmul/matmul-hw.mlir:23273:5
      i_k_next_4028 <= _T_4029;	// matmul/matmul-hw.mlir:23276:7
    else	// matmul/matmul-hw.mlir:23273:5
      i_k_next_4028 <= i_k_next_4025;	// matmul/matmul-hw.mlir:23241:13, :23274:7
  end // always @(posedge)
  assign _T_48 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23278:13
  assign _T_47 = _T_2927 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23279:13
  mult mult_inst247 (	// matmul/matmul-hw.mlir:23280:28
    .a      (A_reg_bank247_p0_rd_data),	// matmul/matmul-hw.mlir:12462:33
    .b      (_T_2581),
    .t      (_T_2927),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst247_result)
  );
  assign _T_46 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23281:13
  assign a_i_k_7_i_j_15 = A_reg_bank247_p0_rd_data;	// matmul/matmul-hw.mlir:12462:33, :23283:5
  //PROBE: a_i_k_7_i_j_15	// matmul/matmul-hw.mlir:23284:5
  assign b_i_k_7_i_j_15 = _T_2581;	// matmul/matmul-hw.mlir:23286:5
  //PROBE: b_i_k_7_i_j_15	// matmul/matmul-hw.mlir:23287:5
  assign c_prev_i_k_7_i_j_15 = C_reg_bank7_p0_rd_data;	// matmul/matmul-hw.mlir:23056:36, :23289:5
  //PROBE: c_prev_i_k_7_i_j_15	// matmul/matmul-hw.mlir:23290:5
  assign tk_i_k_7_i_j_15 = _T_2917;	// matmul/matmul-hw.mlir:23292:5
  //PROBE: tk_i_k_7_i_j_15	// matmul/matmul-hw.mlir:23293:5
  wire [31:0] _T_4030 = mult_inst247_result + C_reg_bank7_p0_rd_data;	// matmul/matmul-hw.mlir:23056:36, :23280:28, :23294:13
  assign c_i_k_7_i_j_15 = _T_4030;	// matmul/matmul-hw.mlir:23296:5
  //PROBE: c_i_k_7_i_j_15	// matmul/matmul-hw.mlir:23297:5
  assign _T_45 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23298:13
  assign _T_44 = _T_2937 ? _T_4030 : 32'bx;	// matmul/matmul-hw.mlir:8079:18, :23299:13
  localparam [3:0] _T_4032 = 4'h0;	// matmul/matmul-hw.mlir:23302:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23303:5
    if (rst)	// matmul/matmul-hw.mlir:23303:5
      i_k_next_4031 <= _T_4032;	// matmul/matmul-hw.mlir:23306:7
    else	// matmul/matmul-hw.mlir:23303:5
      i_k_next_4031 <= i_k_next_4028;	// matmul/matmul-hw.mlir:23271:13, :23304:7
  end // always @(posedge)
  assign _T_43 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23308:13
  assign _T_42 = _T_2932 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23309:13
  mult mult_inst248 (	// matmul/matmul-hw.mlir:23310:28
    .a      (A_reg_bank248_p0_rd_data),	// matmul/matmul-hw.mlir:12463:33
    .b      (_T_2597),
    .t      (_T_2932),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst248_result)
  );
  assign _T_41 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23311:13
  assign a_i_k_8_i_j_15 = A_reg_bank248_p0_rd_data;	// matmul/matmul-hw.mlir:12463:33, :23313:5
  //PROBE: a_i_k_8_i_j_15	// matmul/matmul-hw.mlir:23314:5
  assign b_i_k_8_i_j_15 = _T_2597;	// matmul/matmul-hw.mlir:23316:5
  //PROBE: b_i_k_8_i_j_15	// matmul/matmul-hw.mlir:23317:5
  assign c_prev_i_k_8_i_j_15 = C_reg_bank8_p0_rd_data;	// matmul/matmul-hw.mlir:23057:36, :23319:5
  //PROBE: c_prev_i_k_8_i_j_15	// matmul/matmul-hw.mlir:23320:5
  assign tk_i_k_8_i_j_15 = _T_2922;	// matmul/matmul-hw.mlir:23322:5
  //PROBE: tk_i_k_8_i_j_15	// matmul/matmul-hw.mlir:23323:5
  wire [31:0] _T_4033 = mult_inst248_result + C_reg_bank8_p0_rd_data;	// matmul/matmul-hw.mlir:23057:36, :23310:28, :23324:13
  assign c_i_k_8_i_j_15 = _T_4033;	// matmul/matmul-hw.mlir:23326:5
  //PROBE: c_i_k_8_i_j_15	// matmul/matmul-hw.mlir:23327:5
  assign _T_40 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23328:13
  assign _T_39 = _T_2942 ? _T_4033 : 32'bx;	// matmul/matmul-hw.mlir:8074:18, :23329:13
  localparam [3:0] _T_4035 = 4'h0;	// matmul/matmul-hw.mlir:23332:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23333:5
    if (rst)	// matmul/matmul-hw.mlir:23333:5
      i_k_next_4034 <= _T_4035;	// matmul/matmul-hw.mlir:23336:7
    else	// matmul/matmul-hw.mlir:23333:5
      i_k_next_4034 <= i_k_next_4031;	// matmul/matmul-hw.mlir:23301:13, :23334:7
  end // always @(posedge)
  assign _T_38 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23338:13
  assign _T_37 = _T_2937 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23339:13
  mult mult_inst249 (	// matmul/matmul-hw.mlir:23340:28
    .a      (A_reg_bank249_p0_rd_data),	// matmul/matmul-hw.mlir:12464:33
    .b      (_T_2613),
    .t      (_T_2937),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst249_result)
  );
  assign _T_36 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23341:13
  assign a_i_k_9_i_j_15 = A_reg_bank249_p0_rd_data;	// matmul/matmul-hw.mlir:12464:33, :23343:5
  //PROBE: a_i_k_9_i_j_15	// matmul/matmul-hw.mlir:23344:5
  assign b_i_k_9_i_j_15 = _T_2613;	// matmul/matmul-hw.mlir:23346:5
  //PROBE: b_i_k_9_i_j_15	// matmul/matmul-hw.mlir:23347:5
  assign c_prev_i_k_9_i_j_15 = C_reg_bank9_p0_rd_data;	// matmul/matmul-hw.mlir:23058:36, :23349:5
  //PROBE: c_prev_i_k_9_i_j_15	// matmul/matmul-hw.mlir:23350:5
  assign tk_i_k_9_i_j_15 = _T_2927;	// matmul/matmul-hw.mlir:23352:5
  //PROBE: tk_i_k_9_i_j_15	// matmul/matmul-hw.mlir:23353:5
  wire [31:0] _T_4036 = mult_inst249_result + C_reg_bank9_p0_rd_data;	// matmul/matmul-hw.mlir:23058:36, :23340:28, :23354:13
  assign c_i_k_9_i_j_15 = _T_4036;	// matmul/matmul-hw.mlir:23356:5
  //PROBE: c_i_k_9_i_j_15	// matmul/matmul-hw.mlir:23357:5
  assign _T_35 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23358:13
  assign _T_34 = _T_2947 ? _T_4036 : 32'bx;	// matmul/matmul-hw.mlir:8069:18, :23359:13
  localparam [3:0] _T_4038 = 4'h0;	// matmul/matmul-hw.mlir:23362:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23363:5
    if (rst)	// matmul/matmul-hw.mlir:23363:5
      i_k_next_4037 <= _T_4038;	// matmul/matmul-hw.mlir:23366:7
    else	// matmul/matmul-hw.mlir:23363:5
      i_k_next_4037 <= i_k_next_4034;	// matmul/matmul-hw.mlir:23331:13, :23364:7
  end // always @(posedge)
  assign _T_33 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23368:13
  assign _T_32 = _T_2942 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23369:13
  mult mult_inst250 (	// matmul/matmul-hw.mlir:23370:28
    .a      (A_reg_bank250_p0_rd_data),	// matmul/matmul-hw.mlir:12465:33
    .b      (_T_2629),
    .t      (_T_2942),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst250_result)
  );
  assign _T_31 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23371:13
  assign a_i_k_10_i_j_15 = A_reg_bank250_p0_rd_data;	// matmul/matmul-hw.mlir:12465:33, :23373:5
  //PROBE: a_i_k_10_i_j_15	// matmul/matmul-hw.mlir:23374:5
  assign b_i_k_10_i_j_15 = _T_2629;	// matmul/matmul-hw.mlir:23376:5
  //PROBE: b_i_k_10_i_j_15	// matmul/matmul-hw.mlir:23377:5
  assign c_prev_i_k_10_i_j_15 = C_reg_bank10_p0_rd_data;	// matmul/matmul-hw.mlir:23059:37, :23379:5
  //PROBE: c_prev_i_k_10_i_j_15	// matmul/matmul-hw.mlir:23380:5
  assign tk_i_k_10_i_j_15 = _T_2932;	// matmul/matmul-hw.mlir:23382:5
  //PROBE: tk_i_k_10_i_j_15	// matmul/matmul-hw.mlir:23383:5
  wire [31:0] _T_4039 = mult_inst250_result + C_reg_bank10_p0_rd_data;	// matmul/matmul-hw.mlir:23059:37, :23370:28, :23384:13
  assign c_i_k_10_i_j_15 = _T_4039;	// matmul/matmul-hw.mlir:23386:5
  //PROBE: c_i_k_10_i_j_15	// matmul/matmul-hw.mlir:23387:5
  assign _T_30 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23388:13
  assign _T_29 = _T_2952 ? _T_4039 : 32'bx;	// matmul/matmul-hw.mlir:8064:18, :23389:13
  localparam [3:0] _T_4041 = 4'h0;	// matmul/matmul-hw.mlir:23392:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23393:5
    if (rst)	// matmul/matmul-hw.mlir:23393:5
      i_k_next_4040 <= _T_4041;	// matmul/matmul-hw.mlir:23396:7
    else	// matmul/matmul-hw.mlir:23393:5
      i_k_next_4040 <= i_k_next_4037;	// matmul/matmul-hw.mlir:23361:13, :23394:7
  end // always @(posedge)
  assign _T_28 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23398:13
  assign _T_27 = _T_2947 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23399:13
  mult mult_inst251 (	// matmul/matmul-hw.mlir:23400:28
    .a      (A_reg_bank251_p0_rd_data),	// matmul/matmul-hw.mlir:12466:33
    .b      (_T_2645),
    .t      (_T_2947),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst251_result)
  );
  assign _T_26 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23401:13
  assign a_i_k_11_i_j_15 = A_reg_bank251_p0_rd_data;	// matmul/matmul-hw.mlir:12466:33, :23403:5
  //PROBE: a_i_k_11_i_j_15	// matmul/matmul-hw.mlir:23404:5
  assign b_i_k_11_i_j_15 = _T_2645;	// matmul/matmul-hw.mlir:23406:5
  //PROBE: b_i_k_11_i_j_15	// matmul/matmul-hw.mlir:23407:5
  assign c_prev_i_k_11_i_j_15 = C_reg_bank11_p0_rd_data;	// matmul/matmul-hw.mlir:23060:37, :23409:5
  //PROBE: c_prev_i_k_11_i_j_15	// matmul/matmul-hw.mlir:23410:5
  assign tk_i_k_11_i_j_15 = _T_2937;	// matmul/matmul-hw.mlir:23412:5
  //PROBE: tk_i_k_11_i_j_15	// matmul/matmul-hw.mlir:23413:5
  wire [31:0] _T_4042 = mult_inst251_result + C_reg_bank11_p0_rd_data;	// matmul/matmul-hw.mlir:23060:37, :23400:28, :23414:13
  assign c_i_k_11_i_j_15 = _T_4042;	// matmul/matmul-hw.mlir:23416:5
  //PROBE: c_i_k_11_i_j_15	// matmul/matmul-hw.mlir:23417:5
  assign _T_25 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23418:13
  assign _T_24 = _T_2957 ? _T_4042 : 32'bx;	// matmul/matmul-hw.mlir:8059:18, :23419:13
  localparam [3:0] _T_4044 = 4'h0;	// matmul/matmul-hw.mlir:23422:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23423:5
    if (rst)	// matmul/matmul-hw.mlir:23423:5
      i_k_next_4043 <= _T_4044;	// matmul/matmul-hw.mlir:23426:7
    else	// matmul/matmul-hw.mlir:23423:5
      i_k_next_4043 <= i_k_next_4040;	// matmul/matmul-hw.mlir:23391:13, :23424:7
  end // always @(posedge)
  assign _T_23 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23428:13
  assign _T_22 = _T_2952 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23429:13
  mult mult_inst252 (	// matmul/matmul-hw.mlir:23430:28
    .a      (A_reg_bank252_p0_rd_data),	// matmul/matmul-hw.mlir:12467:33
    .b      (_T_2661),
    .t      (_T_2952),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst252_result)
  );
  assign _T_21 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23431:13
  assign a_i_k_12_i_j_15 = A_reg_bank252_p0_rd_data;	// matmul/matmul-hw.mlir:12467:33, :23433:5
  //PROBE: a_i_k_12_i_j_15	// matmul/matmul-hw.mlir:23434:5
  assign b_i_k_12_i_j_15 = _T_2661;	// matmul/matmul-hw.mlir:23436:5
  //PROBE: b_i_k_12_i_j_15	// matmul/matmul-hw.mlir:23437:5
  assign c_prev_i_k_12_i_j_15 = C_reg_bank12_p0_rd_data;	// matmul/matmul-hw.mlir:23061:37, :23439:5
  //PROBE: c_prev_i_k_12_i_j_15	// matmul/matmul-hw.mlir:23440:5
  assign tk_i_k_12_i_j_15 = _T_2942;	// matmul/matmul-hw.mlir:23442:5
  //PROBE: tk_i_k_12_i_j_15	// matmul/matmul-hw.mlir:23443:5
  wire [31:0] _T_4045 = mult_inst252_result + C_reg_bank12_p0_rd_data;	// matmul/matmul-hw.mlir:23061:37, :23430:28, :23444:13
  assign c_i_k_12_i_j_15 = _T_4045;	// matmul/matmul-hw.mlir:23446:5
  //PROBE: c_i_k_12_i_j_15	// matmul/matmul-hw.mlir:23447:5
  assign _T_20 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23448:13
  assign _T_19 = _T_2962 ? _T_4045 : 32'bx;	// matmul/matmul-hw.mlir:8054:18, :23449:13
  localparam [3:0] _T_4047 = 4'h0;	// matmul/matmul-hw.mlir:23452:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23453:5
    if (rst)	// matmul/matmul-hw.mlir:23453:5
      i_k_next_4046 <= _T_4047;	// matmul/matmul-hw.mlir:23456:7
    else	// matmul/matmul-hw.mlir:23453:5
      i_k_next_4046 <= i_k_next_4043;	// matmul/matmul-hw.mlir:23421:13, :23454:7
  end // always @(posedge)
  assign _T_18 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23458:13
  assign _T_17 = _T_2957 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23459:13
  mult mult_inst253 (	// matmul/matmul-hw.mlir:23460:28
    .a      (A_reg_bank253_p0_rd_data),	// matmul/matmul-hw.mlir:12468:33
    .b      (_T_2677),
    .t      (_T_2957),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst253_result)
  );
  assign _T_16 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23461:13
  assign a_i_k_13_i_j_15 = A_reg_bank253_p0_rd_data;	// matmul/matmul-hw.mlir:12468:33, :23463:5
  //PROBE: a_i_k_13_i_j_15	// matmul/matmul-hw.mlir:23464:5
  assign b_i_k_13_i_j_15 = _T_2677;	// matmul/matmul-hw.mlir:23466:5
  //PROBE: b_i_k_13_i_j_15	// matmul/matmul-hw.mlir:23467:5
  assign c_prev_i_k_13_i_j_15 = C_reg_bank13_p0_rd_data;	// matmul/matmul-hw.mlir:23062:37, :23469:5
  //PROBE: c_prev_i_k_13_i_j_15	// matmul/matmul-hw.mlir:23470:5
  assign tk_i_k_13_i_j_15 = _T_2947;	// matmul/matmul-hw.mlir:23472:5
  //PROBE: tk_i_k_13_i_j_15	// matmul/matmul-hw.mlir:23473:5
  wire [31:0] _T_4048 = mult_inst253_result + C_reg_bank13_p0_rd_data;	// matmul/matmul-hw.mlir:23062:37, :23460:28, :23474:13
  assign c_i_k_13_i_j_15 = _T_4048;	// matmul/matmul-hw.mlir:23476:5
  //PROBE: c_i_k_13_i_j_15	// matmul/matmul-hw.mlir:23477:5
  assign _T_15 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23478:13
  assign _T_14 = _T_3833 ? _T_4048 : 32'bx;	// matmul/matmul-hw.mlir:8049:18, :23479:13
  localparam [3:0] _T_4050 = 4'h0;	// matmul/matmul-hw.mlir:23482:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23483:5
    if (rst)	// matmul/matmul-hw.mlir:23483:5
      i_k_next_4049 <= _T_4050;	// matmul/matmul-hw.mlir:23486:7
    else	// matmul/matmul-hw.mlir:23483:5
      i_k_next_4049 <= i_k_next_4046;	// matmul/matmul-hw.mlir:23451:13, :23484:7
  end // always @(posedge)
  assign _T_13 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23488:13
  assign _T_12 = _T_2962 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23489:13
  mult mult_inst254 (	// matmul/matmul-hw.mlir:23490:28
    .a      (A_reg_bank254_p0_rd_data),	// matmul/matmul-hw.mlir:12469:33
    .b      (_T_2693),
    .t      (_T_2962),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst254_result)
  );
  assign _T_11 = _T_3909 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23491:13
  assign a_i_k_14_i_j_15 = A_reg_bank254_p0_rd_data;	// matmul/matmul-hw.mlir:12469:33, :23493:5
  //PROBE: a_i_k_14_i_j_15	// matmul/matmul-hw.mlir:23494:5
  assign b_i_k_14_i_j_15 = _T_2693;	// matmul/matmul-hw.mlir:23496:5
  //PROBE: b_i_k_14_i_j_15	// matmul/matmul-hw.mlir:23497:5
  assign c_prev_i_k_14_i_j_15 = C_reg_bank14_p0_rd_data;	// matmul/matmul-hw.mlir:23063:37, :23499:5
  //PROBE: c_prev_i_k_14_i_j_15	// matmul/matmul-hw.mlir:23500:5
  assign tk_i_k_14_i_j_15 = _T_2952;	// matmul/matmul-hw.mlir:23502:5
  //PROBE: tk_i_k_14_i_j_15	// matmul/matmul-hw.mlir:23503:5
  wire [31:0] _T_4051 = mult_inst254_result + C_reg_bank14_p0_rd_data;	// matmul/matmul-hw.mlir:23063:37, :23490:28, :23504:13
  assign c_i_k_14_i_j_15 = _T_4051;	// matmul/matmul-hw.mlir:23506:5
  //PROBE: c_i_k_14_i_j_15	// matmul/matmul-hw.mlir:23507:5
  assign _T_10 = _T_3909 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23508:13
  assign _T_9 = _T_3909 ? _T_4051 : 32'bx;	// matmul/matmul-hw.mlir:8044:18, :23509:13
  localparam [3:0] _T_4053 = 4'h0;	// matmul/matmul-hw.mlir:23512:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23513:5
    if (rst)	// matmul/matmul-hw.mlir:23513:5
      i_k_next_4052 <= _T_4053;	// matmul/matmul-hw.mlir:23516:7
    else	// matmul/matmul-hw.mlir:23513:5
      i_k_next_4052 <= i_k_next_4049;	// matmul/matmul-hw.mlir:23481:13, :23514:7
  end // always @(posedge)
  assign _T_8 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23518:13
  assign _T_7 = _T_3833 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23519:13
  mult mult_inst255 (	// matmul/matmul-hw.mlir:23520:28
    .a      (A_reg_bank255_p0_rd_data),	// matmul/matmul-hw.mlir:12470:33
    .b      (_T_2709),
    .t      (_T_3833),
    .clk    (clk),
    .rst    (rst),
    .result (mult_inst255_result)
  );
  assign _T_6 = _T_3985 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23521:13
  assign a_i_k_15_i_j_15 = A_reg_bank255_p0_rd_data;	// matmul/matmul-hw.mlir:12470:33, :23523:5
  //PROBE: a_i_k_15_i_j_15	// matmul/matmul-hw.mlir:23524:5
  assign b_i_k_15_i_j_15 = _T_2709;	// matmul/matmul-hw.mlir:23526:5
  //PROBE: b_i_k_15_i_j_15	// matmul/matmul-hw.mlir:23527:5
  assign c_prev_i_k_15_i_j_15 = C_reg_bank15_p0_rd_data;	// matmul/matmul-hw.mlir:23064:37, :23529:5
  //PROBE: c_prev_i_k_15_i_j_15	// matmul/matmul-hw.mlir:23530:5
  assign tk_i_k_15_i_j_15 = _T_2957;	// matmul/matmul-hw.mlir:23532:5
  //PROBE: tk_i_k_15_i_j_15	// matmul/matmul-hw.mlir:23533:5
  wire [31:0] _T_4054 = mult_inst255_result + C_reg_bank15_p0_rd_data;	// matmul/matmul-hw.mlir:23064:37, :23520:28, :23534:13
  assign c_i_k_15_i_j_15 = _T_4054;	// matmul/matmul-hw.mlir:23536:5
  //PROBE: c_i_k_15_i_j_15	// matmul/matmul-hw.mlir:23537:5
  assign _T_5 = _T_3985 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23538:13
  assign _T_4 = _T_3985 ? _T_4054 : 32'bx;	// matmul/matmul-hw.mlir:8039:18, :23539:13
  localparam [3:0] _T_4056 = 4'h0;	// matmul/matmul-hw.mlir:23542:19
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23543:5
    if (rst)	// matmul/matmul-hw.mlir:23543:5
      i_k_next_4055 <= _T_4056;	// matmul/matmul-hw.mlir:23546:7
    else	// matmul/matmul-hw.mlir:23543:5
      i_k_next_4055 <= i_k_next_4052;	// matmul/matmul-hw.mlir:23511:13, :23544:7
  end // always @(posedge)
  wire [34:0] _T_4058 = _T_4057;	// matmul/matmul-hw.mlir:23549:13
  wire [34:0] _T_4059 = {_T_4058[6'h0+:34], {{_T_2712}}};	// matmul/matmul-hw.mlir:23550:19, :23551:13, :23552:13, :23553:13
  wire [34:0] _T_4060 = {{1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}, {1'h0}};	// matmul/matmul-hw.mlir:23554:19, :23555:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23556:5
    if (rst)	// matmul/matmul-hw.mlir:23556:5
      _T_4057 <= _T_4060;	// matmul/matmul-hw.mlir:23559:7
    else	// matmul/matmul-hw.mlir:23556:5
      _T_4057 <= _T_4059;	// matmul/matmul-hw.mlir:23557:7
  end // always @(posedge)
  wire _T_4061 = _T_4057[6'h22];	// matmul/matmul-hw.mlir:23549:13, :23561:16, :23562:13
  assign _T_3 = _T_4061 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23563:13
  wire [3:0][3:0] _T_4063 = i_delayed_4062;	// matmul/matmul-hw.mlir:23565:13
  wire [3:0][3:0] _T_4064 = {_T_4063[2'h0+:3], {{i_k_next_4055}}};	// matmul/matmul-hw.mlir:23541:13, :23566:19, :23567:13, :23568:13, :23569:13
  wire [3:0][3:0] _T_4065 = {{4'h0}, {4'h0}, {4'h0}, {4'h0}};	// matmul/matmul-hw.mlir:23570:19, :23571:13
  always @(posedge clk) begin	// matmul/matmul-hw.mlir:23572:5
    if (rst)	// matmul/matmul-hw.mlir:23572:5
      i_delayed_4062 <= _T_4065;	// matmul/matmul-hw.mlir:23575:7
    else	// matmul/matmul-hw.mlir:23572:5
      i_delayed_4062 <= _T_4064;	// matmul/matmul-hw.mlir:23573:7
  end // always @(posedge)
  assign _T_2 = _T_4061 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23579:13
  assign _T_1 = _T_4061 ? i_delayed_4062[2'h3] : 4'bx;	// matmul/matmul-hw.mlir:8036:17, :23565:13, :23577:20, :23578:13, :23580:13
  assign _T_0 = _T_4061 ? 1'h1 : 1'h0;	// matmul/matmul-hw.mlir:8029:13, :8033:14, :23581:13
  assign _T = _T_4061 ? C_reg_bank16_p0_rd_data : 32'bx;	// matmul/matmul-hw.mlir:8034:18, :23065:37, :23582:13
  assign A_p0_addr_en = {{_T_2115}, {_T_2120}, {_T_2125}, {_T_2130}, {_T_2135}, {_T_2140}, {_T_2145}, {_T_2150}, {_T_2155}, {_T_2160}, {_T_2165}, {_T_2170}, {_T_2175}, {_T_2180}, {_T_2185}, {_T_2192}};	// matmul/matmul-hw.mlir:7668:10, :12472:12, :12504:12, :12550:12, :12596:12, :12642:12, :12688:12, :12734:12, :12780:12, :12826:12, :12872:12, :12918:12, :12964:12, :13010:12, :13056:12, :13102:12, :13148:12, :23583:5
  assign A_p0_addr_data = {{_T_2114}, {_T_2119}, {_T_2124}, {_T_2129}, {_T_2134}, {_T_2139}, {_T_2144}, {_T_2149}, {_T_2154}, {_T_2159}, {_T_2164}, {_T_2169}, {_T_2174}, {_T_2179}, {_T_2184}, {_T_2191}};	// matmul/matmul-hw.mlir:7685:10, :12473:12, :12505:12, :12551:12, :12597:12, :12643:12, :12689:12, :12735:12, :12781:12, :12827:12, :12873:12, :12919:12, :12965:12, :13011:12, :13057:12, :13103:12, :13149:12, :23583:5
  assign A_p0_rd_en = {{_T_2113}, {_T_2118}, {_T_2123}, {_T_2128}, {_T_2133}, {_T_2138}, {_T_2143}, {_T_2148}, {_T_2153}, {_T_2158}, {_T_2163}, {_T_2168}, {_T_2173}, {_T_2178}, {_T_2183}, {_T_2190}};	// matmul/matmul-hw.mlir:7702:10, :12474:12, :12506:12, :12552:12, :12598:12, :12644:12, :12690:12, :12736:12, :12782:12, :12828:12, :12874:12, :12920:12, :12966:12, :13012:12, :13058:12, :13104:12, :13150:12, :23583:5
  assign B_p0_rd_en = {{_T_7}, {_T_94}, {_T_181}, {_T_268}, {_T_355}, {_T_442}, {_T_529}, {_T_616}, {_T_703}, {_T_790}, {_T_877}, {_T_964}, {_T_1051}, {_T_1138}, {_T_1225}, {_T_1312}, {_T_12}, {_T_99}, {_T_186}, {_T_273}, {_T_360}, {_T_447}, {_T_534}, {_T_621}, {_T_708}, {_T_795}, {_T_882}, {_T_969}, {_T_1056}, {_T_1143}, {_T_1230}, {_T_1317}, {_T_17}, {_T_104}, {_T_191}, {_T_278}, {_T_365}, {_T_452}, {_T_539}, {_T_626}, {_T_713}, {_T_800}, {_T_887}, {_T_974}, {_T_1061}, {_T_1148}, {_T_1235}, {_T_1322}, {_T_22}, {_T_109}, {_T_196}, {_T_283}, {_T_370}, {_T_457}, {_T_544}, {_T_631}, {_T_718}, {_T_805}, {_T_892}, {_T_979}, {_T_1066}, {_T_1153}, {_T_1240}, {_T_1327}, {_T_27}, {_T_114}, {_T_201}, {_T_288}, {_T_375}, {_T_462}, {_T_549}, {_T_636}, {_T_723}, {_T_810}, {_T_897}, {_T_984}, {_T_1071}, {_T_1158}, {_T_1245}, {_T_1332}, {_T_32}, {_T_119}, {_T_206}, {_T_293}, {_T_380}, {_T_467}, {_T_554}, {_T_641}, {_T_728}, {_T_815}, {_T_902}, {_T_989}, {_T_1076}, {_T_1163}, {_T_1250}, {_T_1337}, {_T_37}, {_T_124}, {_T_211}, {_T_298}, {_T_385}, {_T_472}, {_T_559}, {_T_646}, {_T_733}, {_T_820}, {_T_907}, {_T_994}, {_T_1081}, {_T_1168}, {_T_1255}, {_T_1342}, {_T_42}, {_T_129}, {_T_216}, {_T_303}, {_T_390}, {_T_477}, {_T_564}, {_T_651}, {_T_738}, {_T_825}, {_T_912}, {_T_999}, {_T_1086}, {_T_1173}, {_T_1260}, {_T_1347}, {_T_47}, {_T_134}, {_T_221}, {_T_308}, {_T_395}, {_T_482}, {_T_569}, {_T_656}, {_T_743}, {_T_830}, {_T_917}, {_T_1004}, {_T_1091}, {_T_1178}, {_T_1265}, {_T_1352}, {_T_52}, {_T_139}, {_T_226}, {_T_313}, {_T_400}, {_T_487}, {_T_574}, {_T_661}, {_T_748}, {_T_835}, {_T_922}, {_T_1009}, {_T_1096}, {_T_1183}, {_T_1270}, {_T_1357}, {_T_57}, {_T_144}, {_T_231}, {_T_318}, {_T_405}, {_T_492}, {_T_579}, {_T_666}, {_T_753}, {_T_840}, {_T_927}, {_T_1014}, {_T_1101}, {_T_1188}, {_T_1275}, {_T_1362}, {_T_62}, {_T_149}, {_T_236}, {_T_323}, {_T_410}, {_T_497}, {_T_584}, {_T_671}, {_T_758}, {_T_845}, {_T_932}, {_T_1019}, {_T_1106}, {_T_1193}, {_T_1280}, {_T_1367}, {_T_67}, {_T_154}, {_T_241}, {_T_328}, {_T_415}, {_T_502}, {_T_589}, {_T_676}, {_T_763}, {_T_850}, {_T_937}, {_T_1024}, {_T_1111}, {_T_1198}, {_T_1285}, {_T_1372}, {_T_72}, {_T_159}, {_T_246}, {_T_333}, {_T_420}, {_T_507}, {_T_594}, {_T_681}, {_T_768}, {_T_855}, {_T_942}, {_T_1029}, {_T_1116}, {_T_1203}, {_T_1290}, {_T_1377}, {_T_77}, {_T_164}, {_T_251}, {_T_338}, {_T_425}, {_T_512}, {_T_599}, {_T_686}, {_T_773}, {_T_860}, {_T_947}, {_T_1034}, {_T_1121}, {_T_1208}, {_T_1295}, {_T_1382}, {_T_82}, {_T_169}, {_T_256}, {_T_343}, {_T_430}, {_T_517}, {_T_604}, {_T_691}, {_T_778}, {_T_865}, {_T_952}, {_T_1039}, {_T_1126}, {_T_1213}, {_T_1300}, {_T_1387}};	// matmul/matmul-hw.mlir:7959:10, :14227:13, :14249:13, :14271:13, :14293:13, :14315:13, :14337:13, :14359:13, :14381:13, :14403:13, :14425:13, :14447:13, :14469:13, :14491:13, :14513:13, :14535:13, :14557:13, :14694:13, :14724:13, :14754:13, :14784:13, :14814:13, :14844:13, :14874:13, :14904:13, :14934:13, :14964:13, :14994:13, :15024:13, :15054:13, :15084:13, :15114:13, :15144:13, :15289:13, :15319:13, :15349:13, :15379:13, :15409:13, :15439:13, :15469:13, :15499:13, :15529:13, :15559:13, :15589:13, :15619:13, :15649:13, :15679:13, :15709:13, :15739:13, :15884:13, :15914:13, :15944:13, :15974:13, :16004:13, :16034:13, :16064:13, :16094:13, :16124:13, :16154:13, :16184:13, :16214:13, :16244:13, :16274:13, :16304:13, :16334:13, :16479:13, :16509:13, :16539:13, :16569:13, :16599:13, :16629:13, :16659:13, :16689:13, :16719:13, :16749:13, :16779:13, :16809:13, :16839:13, :16869:13, :16899:13, :16929:13, :17074:13, :17104:13, :17134:13, :17164:13, :17194:13, :17224:13, :17254:13, :17284:13, :17314:13, :17344:13, :17374:13, :17404:13, :17434:13, :17464:13, :17494:13, :17524:13, :17669:13, :17699:13, :17729:13, :17759:13, :17789:13, :17819:13, :17849:13, :17879:13, :17909:13, :17939:13, :17969:13, :17999:13, :18029:13, :18059:13, :18089:13, :18119:13, :18264:13, :18294:13, :18324:13, :18354:13, :18384:13, :18414:13, :18444:13, :18474:13, :18504:13, :18534:13, :18564:13, :18594:13, :18624:13, :18654:13, :18684:13, :18714:13, :18859:13, :18889:13, :18919:13, :18949:13, :18979:13, :19009:13, :19039:13, :19069:13, :19099:13, :19129:13, :19159:13, :19189:13, :19219:13, :19249:13, :19279:13, :19309:13, :19454:13, :19484:13, :19514:13, :19544:13, :19574:13, :19604:13, :19634:13, :19664:13, :19694:13, :19724:13, :19754:13, :19784:13, :19814:13, :19844:13, :19874:13, :19904:13, :20049:13, :20079:13, :20109:13, :20139:13, :20169:13, :20199:13, :20229:13, :20259:13, :20289:13, :20319:13, :20349:13, :20379:13, :20409:13, :20439:13, :20469:13, :20499:13, :20644:13, :20674:13, :20704:13, :20734:13, :20764:13, :20794:13, :20824:13, :20854:13, :20884:13, :20914:13, :20944:13, :20974:13, :21004:13, :21034:13, :21064:13, :21094:13, :21239:13, :21269:13, :21299:13, :21329:13, :21359:13, :21389:13, :21419:13, :21449:13, :21479:13, :21509:13, :21539:13, :21569:13, :21599:13, :21629:13, :21659:13, :21689:13, :21849:13, :21879:13, :21909:13, :21939:13, :21969:13, :21999:13, :22029:13, :22059:13, :22089:13, :22119:13, :22149:13, :22179:13, :22209:13, :22239:13, :22269:13, :22299:13, :22459:13, :22489:13, :22519:13, :22549:13, :22579:13, :22609:13, :22639:13, :22669:13, :22699:13, :22729:13, :22759:13, :22789:13, :22819:13, :22849:13, :22879:13, :22909:13, :23069:13, :23099:13, :23129:13, :23159:13, :23189:13, :23219:13, :23249:13, :23279:13, :23309:13, :23339:13, :23369:13, :23399:13, :23429:13, :23459:13, :23489:13, :23519:13, :23583:5
  assign C_p0_addr_en = {{_T_2}, {_T_89}, {_T_176}, {_T_263}, {_T_350}, {_T_437}, {_T_524}, {_T_611}, {_T_698}, {_T_785}, {_T_872}, {_T_959}, {_T_1046}, {_T_1133}, {_T_1220}, {_T_1307}};	// matmul/matmul-hw.mlir:7976:10, :14594:13, :15189:13, :15784:13, :16379:13, :16974:13, :17569:13, :18164:13, :18759:13, :19354:13, :19949:13, :20544:13, :21139:13, :21749:13, :22359:13, :22969:13, :23579:13, :23583:5
  assign C_p0_addr_data = {{_T_1}, {_T_88}, {_T_175}, {_T_262}, {_T_349}, {_T_436}, {_T_523}, {_T_610}, {_T_697}, {_T_784}, {_T_871}, {_T_958}, {_T_1045}, {_T_1132}, {_T_1219}, {_T_1306}};	// matmul/matmul-hw.mlir:7993:10, :14595:13, :15190:13, :15785:13, :16380:13, :16975:13, :17570:13, :18165:13, :18760:13, :19355:13, :19950:13, :20545:13, :21140:13, :21750:13, :22360:13, :22970:13, :23580:13, :23583:5
  assign C_p0_wr_en = {{_T_0}, {_T_87}, {_T_174}, {_T_261}, {_T_348}, {_T_435}, {_T_522}, {_T_609}, {_T_696}, {_T_783}, {_T_870}, {_T_957}, {_T_1044}, {_T_1131}, {_T_1218}, {_T_1305}};	// matmul/matmul-hw.mlir:8010:10, :14596:13, :15191:13, :15786:13, :16381:13, :16976:13, :17571:13, :18166:13, :18761:13, :19356:13, :19951:13, :20546:13, :21141:13, :21751:13, :22361:13, :22971:13, :23581:13, :23583:5
  assign C_p0_wr_data = {{_T}, {_T_86}, {_T_173}, {_T_260}, {_T_347}, {_T_434}, {_T_521}, {_T_608}, {_T_695}, {_T_782}, {_T_869}, {_T_956}, {_T_1043}, {_T_1130}, {_T_1217}, {_T_1304}};	// matmul/matmul-hw.mlir:8027:10, :14597:13, :15192:13, :15787:13, :16382:13, :16977:13, :17572:13, :18167:13, :18762:13, :19357:13, :19952:13, :20547:13, :21142:13, :21752:13, :22362:13, :22972:13, :23582:13, :23583:5
endmodule

